/home/aavyas1/research/Jonti_Transfers/SLM_RAS/FP_Units/apr_16/mult_16/asap7_tech_4x_170803.lef