/home/aavyas1/research/Jonti_Transfers/SLM_RAS/FP_Units/apr_32/adder32/asap7_tech_4x_170803.lef