/home/aavyas1/research/Jonti_Transfers/SLM_RAS/FP_Units/apr_32/adder32/asap7sc7p5t_24_R_4x_170912.lef