VERSION 5.8 ; 
BUSBITCHARS "[]" ; 
DIVIDERCHAR "/" ; 

PROPERTYDEFINITIONS 
MACRO oaTaper STRING ; 
END PROPERTYDEFINITIONS 

MACRO A2O1A1Ixp33_ASAP7_75t_R_v1 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN A2O1A1Ixp33_ASAP7_75t_R_v1 0 0 ; 
SIZE 1.728 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.224 0.432 0.296 0.936 ; 
RECT 0.088 0.864 0.296 0.936 ; 
RECT 0.224 0.432 0.396 0.504 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.432 0.576 0.816 ; 
RECT 0.504 0.432 0.684 0.504 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.36 1.008 0.7 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.152 0.288 1.224 0.7 ; 
RECT 1.152 0.288 1.324 0.36 ; 
END 
END C 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.304 0.144 1.544 0.216 ; 
RECT 1.472 0.144 1.544 0.936 ; 
RECT 1.024 0.864 1.544 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.728 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.728 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.072 0.252 0.856 0.324 ; 
RECT 0.072 0.252 0.144 0.74 ; 
RECT 0.784 0.252 0.856 0.924 ; 
RECT 0.16 0.108 1.136 0.18 ; 
END 
END A2O1A1Ixp33_ASAP7_75t_R_v1 

MACRO A2O1A1Ixp33_ASAP7_75t_R_v2 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN A2O1A1Ixp33_ASAP7_75t_R_v2 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.152 0.288 0.336 0.36 ; 
RECT 0.264 0.288 0.336 0.792 ; 
RECT 0.192 0.72 0.416 0.792 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.288 0.576 0.668 ; 
RECT 0.504 0.288 0.672 0.36 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.432 0.792 0.668 ; 
RECT 0.824 0.292 0.896 0.504 ; 
RECT 0.72 0.432 0.896 0.504 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.024 0.288 1.224 0.36 ; 
RECT 1.152 0.288 1.224 0.668 ; 
END 
END C 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.216 0.144 1.44 0.216 ; 
RECT 1.368 0.144 1.44 0.936 ; 
RECT 1 0.864 1.44 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 0.704 0.972 ; 
RECT 0.16 0.108 0.916 0.18 ; 
END 
END A2O1A1Ixp33_ASAP7_75t_R_v2 

MACRO A2O1A1O1Ixp33_ASAP7_75t_R_v1 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN A2O1A1O1Ixp33_ASAP7_75t_R_v1 0 0 ; 
SIZE 1.944 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.464 0.576 0.648 ; 
RECT 0.412 0.576 0.576 0.648 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.484 0.792 0.648 ; 
RECT 0.988 0.288 1.06 0.648 ; 
RECT 0.72 0.576 1.06 0.648 ; 
RECT 0.988 0.288 1.144 0.36 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.124 0.432 0.292 0.504 ; 
RECT 0.22 0.432 0.292 0.596 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.284 0.288 1.448 0.36 ; 
RECT 1.376 0.288 1.448 0.648 ; 
RECT 1.228 0.576 1.448 0.648 ; 
END 
END C 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.56 0.288 1.724 0.36 ; 
RECT 1.652 0.288 1.724 0.936 ; 
RECT 1.652 0.864 1.82 0.936 ; 
END 
END D 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.144 1.876 0.216 ; 
RECT 1.804 0.144 1.876 0.672 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.944 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.944 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.18 0.16 0.252 0.36 ; 
RECT 0.18 0.288 0.888 0.36 ; 
RECT 0.38 0.9 0.92 0.972 ; 
RECT 0.184 0.756 1.548 0.828 ; 
RECT 0.184 0.756 0.256 0.936 ; 
RECT 1.476 0.756 1.548 0.944 ; 
END 
END A2O1A1O1Ixp33_ASAP7_75t_R_v1 

MACRO A2O1A1O1Ixp33_ASAP7_75t_R_v2 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN A2O1A1O1Ixp33_ASAP7_75t_R_v2 0 0 ; 
SIZE 1.944 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.288 0.576 0.792 ; 
RECT 0.412 0.72 0.576 0.792 ; 
RECT 0.504 0.288 0.676 0.36 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.108 0.288 0.288 0.36 ; 
RECT 0.216 0.288 0.288 0.668 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.724 0.492 0.796 0.668 ; 
END 
END C 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.94 0.288 1.012 0.668 ; 
RECT 0.94 0.288 1.148 0.36 ; 
END 
END D 
PIN E 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.368 0.288 1.44 0.792 ; 
RECT 1.244 0.72 1.44 0.792 ; 
RECT 1.368 0.288 1.544 0.36 ; 
RECT 1.156 0.508 1.656 0.58 ; 
END 
END E 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.036 0.108 1.872 0.18 ; 
RECT 1.8 0.108 1.872 0.796 ; 
RECT 1.692 0.724 1.872 0.796 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.944 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.944 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 0.704 0.972 ; 
RECT 0.16 0.108 0.908 0.18 ; 
RECT 0.828 0.776 0.9 0.972 ; 
RECT 0.828 0.9 1.568 0.972 ; 
END 
END A2O1A1O1Ixp33_ASAP7_75t_R_v2 

MACRO A2O1Ixp5_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN A2O1Ixp5_ASAP7_75t_R 0 0 ; 
SIZE 1.08 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.412 0.576 0.792 ; 
RECT 0.384 0.72 0.576 0.792 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.16 0.36 0.6 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.316 0.792 0.608 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.592 0.144 1.008 0.216 ; 
RECT 0.936 0.144 1.008 0.84 ; 
RECT 0.804 0.768 1.008 0.84 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.08 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.08 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 0.704 0.972 ; 
END 
END A2O1Ixp5_ASAP7_75t_R 

MACRO AND4x2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AND4x2_ASAP7_75t_R 0 0 ; 
SIZE 3.456 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.12 0.288 0.292 0.36 ; 
RECT 0.22 0.288 0.292 0.792 ; 
RECT 0.104 0.72 0.292 0.792 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.876 0.432 1.036 0.504 ; 
RECT 0.964 0.432 1.036 0.792 ; 
RECT 0.848 0.72 1.036 0.792 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.38 0.432 1.62 0.504 ; 
RECT 1.548 0.432 1.62 0.792 ; 
RECT 1.548 0.72 1.712 0.792 ; 
END 
END C 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.268 0.288 2.34 0.648 ; 
RECT 2.164 0.576 2.34 0.648 ; 
RECT 2.268 0.288 2.48 0.36 ; 
END 
END D 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.972 0.144 3.396 0.216 ; 
RECT 3.324 0.144 3.396 0.936 ; 
RECT 2.972 0.864 3.396 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.456 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.456 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.164 0.116 1.128 0.188 ; 
RECT 0.812 0.284 1.784 0.356 ; 
RECT 1.456 0.116 2.424 0.188 ; 
RECT 0.396 0.336 0.468 0.716 ; 
RECT 0.396 0.644 0.576 0.716 ; 
RECT 2.84 0.448 2.912 0.8 ; 
RECT 2.448 0.728 2.912 0.8 ; 
RECT 0.504 0.644 0.576 0.972 ; 
RECT 2.448 0.728 2.52 0.972 ; 
RECT 0.376 0.9 2.52 0.972 ; 
END 
END AND4x2_ASAP7_75t_R 

MACRO AO21x2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AO21x2_ASAP7_75t_R 0 0 ; 
SIZE 1.944 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.408 0.36 0.656 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.412 0.576 0.656 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.412 0.792 0.656 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.24 0.144 1.868 0.216 ; 
RECT 1.796 0.144 1.868 0.936 ; 
RECT 1.24 0.864 1.868 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.944 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.944 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 0.704 0.972 ; 
RECT 0.16 0.108 1.008 0.18 ; 
RECT 0.936 0.5 1.676 0.572 ; 
RECT 0.936 0.108 1.008 0.828 ; 
RECT 0.696 0.756 1.008 0.828 ; 
END 
END AO21x2_ASAP7_75t_R 

MACRO AO22x2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AO22x2_ASAP7_75t_R 0 0 ; 
SIZE 2.16 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.116 0.504 0.188 0.668 ; 
RECT 0.116 0.504 0.38 0.576 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.482 0.576 0.792 ; 
RECT 0.34 0.72 0.576 0.792 ; 
END 
END A2 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.288 1.008 0.596 ; 
RECT 0.936 0.288 1.148 0.36 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.412 0.792 0.596 ; 
END 
END B2 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.672 0.144 2.092 0.216 ; 
RECT 2.02 0.144 2.092 0.936 ; 
RECT 1.672 0.864 2.092 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.16 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.16 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 1.136 0.972 ; 
RECT 0.592 0.108 1.404 0.18 ; 
RECT 1.332 0.5 1.676 0.572 ; 
RECT 1.332 0.108 1.404 0.828 ; 
RECT 0.808 0.756 1.404 0.828 ; 
END 
END AO22x2_ASAP7_75t_R 

MACRO AO31x2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AO31x2_ASAP7_75t_R 0 0 ; 
SIZE 3.456 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.536 0.268 2.608 0.576 ; 
RECT 2.2 0.504 2.608 0.576 ; 
RECT 2.536 0.268 2.692 0.34 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.268 0.412 1.432 0.484 ; 
RECT 1.36 0.412 1.432 0.576 ; 
RECT 1.36 0.504 1.712 0.576 ; 
RECT 1.64 0.504 1.712 0.668 ; 
RECT 1.64 0.596 1.796 0.668 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.196 0.268 0.36 0.34 ; 
RECT 0.288 0.268 0.36 0.812 ; 
RECT 0.196 0.74 0.36 0.812 ; 
END 
END A3 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.624 0.284 0.696 0.8 ; 
RECT 0.624 0.504 0.792 0.576 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.968 0.108 3.384 0.18 ; 
RECT 3.312 0.108 3.384 0.972 ; 
RECT 2.964 0.9 3.384 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.456 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.456 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.384 0.108 1.788 0.18 ; 
RECT 0.164 0.9 2.216 0.972 ; 
RECT 1.472 0.252 2.424 0.324 ; 
RECT 2.104 0.108 2.864 0.18 ; 
RECT 0.8 0.252 1.104 0.324 ; 
RECT 2.792 0.504 3.188 0.576 ; 
RECT 1.032 0.252 1.104 0.812 ; 
RECT 0.796 0.74 2.42 0.812 ; 
RECT 2.348 0.74 2.42 0.972 ; 
RECT 2.792 0.108 2.864 0.972 ; 
RECT 2.348 0.9 2.864 0.972 ; 
END 
END AO31x2_ASAP7_75t_R 

MACRO AO32x2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AO32x2_ASAP7_75t_R 0 0 ; 
SIZE 2.376 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.132 0.252 0.292 0.324 ; 
RECT 0.22 0.252 0.292 0.972 ; 
RECT 0.132 0.9 0.292 0.972 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.416 0.252 0.576 0.324 ; 
RECT 0.504 0.252 0.576 0.812 ; 
RECT 0.416 0.728 0.576 0.812 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.408 0.792 0.812 ; 
RECT 0.72 0.74 0.888 0.812 ; 
END 
END A3 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.268 1.008 0.608 ; 
RECT 0.936 0.268 1.104 0.34 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.22 0.268 1.292 0.668 ; 
RECT 1.22 0.268 1.408 0.34 ; 
RECT 1.22 0.596 1.42 0.668 ; 
END 
END B2 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.888 0.108 2.088 0.18 ; 
RECT 2.016 0.108 2.088 0.972 ; 
RECT 1.888 0.9 2.088 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.376 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.376 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.392 0.9 1.352 0.972 ; 
RECT 0.16 0.108 1.656 0.18 ; 
RECT 1.584 0.508 1.84 0.58 ; 
RECT 1.584 0.108 1.656 0.828 ; 
RECT 1.04 0.756 1.656 0.828 ; 
END 
END AO32x2_ASAP7_75t_R 

MACRO AOI211xp5_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI211xp5_ASAP7_75t_R 0 0 ; 
SIZE 2.808 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.736 0.252 0.896 0.324 ; 
RECT 0.824 0.252 0.896 0.828 ; 
RECT 0.724 0.756 0.896 0.828 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.312 0.252 0.472 0.324 ; 
RECT 0.4 0.252 0.472 0.828 ; 
RECT 0.3 0.756 0.472 0.828 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.584 0.252 1.656 0.684 ; 
RECT 1.584 0.252 1.768 0.324 ; 
RECT 1.584 0.612 1.768 0.684 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.012 0.252 2.196 0.324 ; 
RECT 2.124 0.252 2.196 0.684 ; 
RECT 2.012 0.612 2.196 0.684 ; 
END 
END C 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.316 0.504 2.388 0.828 ; 
RECT 2.076 0.756 2.388 0.828 ; 
RECT 0.364 0.108 2.524 0.18 ; 
RECT 2.452 0.108 2.524 0.576 ; 
RECT 2.316 0.504 2.524 0.576 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.808 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.808 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 1.152 0.756 1.796 0.828 ; 
RECT 1.152 0.756 1.224 0.972 ; 
RECT 0.364 0.9 1.224 0.972 ; 
RECT 1.444 0.9 2.432 0.972 ; 
END 
END AOI211xp5_ASAP7_75t_R 

MACRO AOI21_x2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI21_x2_ASAP7_75t_R 0 0 ; 
SIZE 1.08 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.184 0.268 0.36 0.34 ; 
RECT 0.288 0.268 0.36 0.812 ; 
RECT 0.188 0.74 0.36 0.812 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.264 0.576 0.656 ; 
RECT 0.504 0.264 0.68 0.336 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.412 0.792 0.812 ; 
RECT 0.62 0.74 0.792 0.812 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.16 0.108 1.008 0.18 ; 
RECT 0.936 0.108 1.008 0.972 ; 
RECT 0.82 0.9 1.008 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.08 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.08 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 0.688 0.972 ; 
END 
END AOI21_x2_ASAP7_75t_R 

MACRO AOI221xp5_ASAP_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI221xp5_ASAP_75t_R 0 0 ; 
SIZE 3.024 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.724 0.108 0.892 0.18 ; 
RECT 0.82 0.108 0.892 0.576 ; 
RECT 0.716 0.504 1.012 0.576 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.272 0.108 0.46 0.18 ; 
RECT 0.388 0.108 0.46 0.576 ; 
RECT 0.284 0.504 0.58 0.576 ; 
END 
END A2 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.128 0.324 1.328 0.396 ; 
RECT 1.256 0.324 1.328 0.576 ; 
RECT 1.256 0.504 1.444 0.576 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2 0.324 2.168 0.396 ; 
RECT 1.788 0.504 2.168 0.576 ; 
RECT 2.096 0.324 2.168 0.828 ; 
RECT 2.096 0.756 2.26 0.828 ; 
END 
END B2 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.268 0.324 2.436 0.396 ; 
RECT 2.36 0.324 2.432 0.8 ; 
RECT 2.36 0.324 2.436 0.576 ; 
RECT 2.36 0.504 2.536 0.576 ; 
END 
END C 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.032 0.18 2.95 0.252 ; 
RECT 2.878 0.18 2.95 0.828 ; 
RECT 2.544 0.756 2.95 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.024 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.024 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.168 0.72 1.992 0.792 ; 
RECT 1.248 0.9 2.856 0.972 ; 
END 
END AOI221xp5_ASAP_75t_R 

MACRO AOI22xp33_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI22xp33_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.116 0.504 0.188 0.668 ; 
RECT 0.116 0.504 0.38 0.576 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.482 0.576 0.792 ; 
RECT 0.34 0.72 0.576 0.792 ; 
END 
END A2 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.924 0.252 1.076 0.324 ; 
RECT 1.004 0.252 1.076 0.596 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.412 0.792 0.596 ; 
END 
END B2 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.592 0.108 1.224 0.18 ; 
RECT 1.152 0.108 1.224 0.828 ; 
RECT 0.808 0.756 1.224 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 1.136 0.972 ; 
END 
END AOI22xp33_ASAP7_75t_R 

MACRO AOI31xp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI31xp67_ASAP7_75t_R 0 0 ; 
SIZE 2.808 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.524 0.288 2.596 0.576 ; 
RECT 2.2 0.504 2.596 0.576 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.288 0.288 1.36 0.576 ; 
RECT 1.288 0.504 1.712 0.576 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.196 0.272 0.36 0.344 ; 
RECT 0.288 0.272 0.36 0.816 ; 
RECT 0.196 0.744 0.36 0.816 ; 
END 
END A3 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.624 0.28 0.696 0.796 ; 
RECT 0.624 0.504 0.852 0.576 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.104 0.108 2.688 0.18 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.808 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.808 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.384 0.108 1.788 0.18 ; 
RECT 0.164 0.9 2.216 0.972 ; 
RECT 1.464 0.312 2.424 0.384 ; 
RECT 0.8 0.252 1.112 0.324 ; 
RECT 1.04 0.252 1.112 0.808 ; 
RECT 0.796 0.736 2.688 0.808 ; 
END 
END AOI31xp67_ASAP7_75t_R 

MACRO AOI322xp5_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI322xp5_ASAP7_75t_R 0 0 ; 
SIZE 2.376 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.116 0.252 0.292 0.324 ; 
RECT 0.22 0.252 0.292 0.604 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.412 0.252 0.576 0.324 ; 
RECT 0.504 0.252 0.576 0.656 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.28 0.792 0.656 ; 
END 
END A3 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.22 0.252 1.292 0.656 ; 
RECT 1.22 0.252 1.384 0.324 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.252 1.008 0.656 ; 
RECT 0.936 0.252 1.1 0.324 ; 
END 
END B2 
PIN C1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.708 0.252 1.872 0.324 ; 
RECT 1.8 0.252 1.872 0.656 ; 
END 
END C1 
PIN C2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.016 0.136 2.088 0.656 ; 
END 
END C2 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.484 0.108 1.556 0.828 ; 
RECT 0.168 0.108 1.776 0.18 ; 
RECT 2.236 0.176 2.308 0.828 ; 
RECT 1.484 0.756 2.308 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.376 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.376 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.384 0.756 1.344 0.828 ; 
RECT 1.032 0.9 1.992 0.972 ; 
END 
END AOI322xp5_ASAP7_75t_R 

MACRO AOI32xp33_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI32xp33_ASAP7_75t_R 0 0 ; 
SIZE 1.728 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.132 0.252 0.292 0.324 ; 
RECT 0.22 0.252 0.292 0.972 ; 
RECT 0.132 0.9 0.292 0.972 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.416 0.252 0.576 0.324 ; 
RECT 0.504 0.252 0.576 0.812 ; 
RECT 0.416 0.728 0.576 0.812 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.408 0.792 0.812 ; 
RECT 0.72 0.74 0.888 0.812 ; 
END 
END A3 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.268 1.008 0.608 ; 
RECT 0.936 0.268 1.104 0.34 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.22 0.268 1.292 0.668 ; 
RECT 1.22 0.268 1.408 0.34 ; 
RECT 1.22 0.596 1.42 0.668 ; 
END 
END B2 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.16 0.108 1.604 0.18 ; 
RECT 1.532 0.108 1.604 0.828 ; 
RECT 1.04 0.756 1.604 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.728 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.728 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.392 0.9 1.336 0.972 ; 
END 
END AOI32xp33_ASAP7_75t_R 

MACRO AOI333xp33_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI333xp33_ASAP7_75t_R 0 0 ; 
SIZE 2.376 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.28 0.792 0.656 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.28 0.576 0.656 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.28 0.36 0.656 ; 
END 
END A3 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.28 1.008 0.656 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.152 0.28 1.224 0.656 ; 
END 
END B2 
PIN B3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.368 0.28 1.44 0.656 ; 
END 
END B3 
PIN C1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.016 0.28 2.088 0.8 ; 
END 
END C1 
PIN C2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.8 0.28 1.872 0.8 ; 
END 
END C2 
PIN C3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.584 0.28 1.656 0.8 ; 
END 
END C3 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.084 0.108 0.156 0.972 ; 
RECT 0.084 0.9 0.732 0.972 ; 
RECT 0.084 0.108 2.27 0.18 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.376 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.376 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.308 0.756 1.4 0.828 ; 
RECT 0.968 0.9 2.06 0.972 ; 
END 
END AOI333xp33_ASAP7_75t_R 

MACRO AOI33xp33_ASAP_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN AOI33xp33_ASAP_75t_R 0 0 ; 
SIZE 1.944 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.068 0.108 0.14 0.576 ; 
RECT 0.068 0.108 0.252 0.18 ; 
RECT 0.288 0.412 0.36 0.576 ; 
RECT 0.068 0.504 0.36 0.576 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.068 0.648 0.14 0.972 ; 
RECT 0.068 0.9 0.244 0.972 ; 
RECT 0.504 0.408 0.576 0.72 ; 
RECT 0.068 0.648 0.576 0.72 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.48 0.792 0.828 ; 
RECT 0.72 0.756 0.892 0.828 ; 
END 
END A3 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.832 0.268 1.008 0.344 ; 
RECT 0.936 0.268 1.008 0.564 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.152 0.268 1.224 0.58 ; 
RECT 1.152 0.268 1.328 0.34 ; 
END 
END B2 
PIN B3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.436 0.412 1.508 0.68 ; 
RECT 1.436 0.412 1.608 0.484 ; 
RECT 1.436 0.608 1.608 0.68 ; 
END 
END B3 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.804 0.108 1.872 0.18 ; 
RECT 1.8 0.108 1.872 0.828 ; 
RECT 1.024 0.756 1.872 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.944 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.944 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.388 0.9 1.352 0.972 ; 
END 
END AOI33xp33_ASAP_75t_R 

MACRO BUFx10_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN BUFx10_ASAP7_75t_R 0 0 ; 
SIZE 3.456 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.288 0.292 0.792 ; 
RECT 0.12 0.72 0.292 0.792 ; 
RECT 0.22 0.288 0.384 0.36 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.024 0.144 3.388 0.216 ; 
RECT 3.316 0.144 3.388 0.936 ; 
RECT 1.022 0.864 3.388 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.456 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.456 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.108 0.796 0.18 ; 
RECT 0.724 0.504 3.186 0.576 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.16 0.9 0.796 0.972 ; 
END 
END BUFx10_ASAP7_75t_R 

MACRO BUFx12_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN BUFx12_ASAP7_75t_R 0 0 ; 
SIZE 3.888 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.24 0.144 3.816 0.216 ; 
RECT 3.744 0.144 3.816 0.936 ; 
RECT 1.24 0.864 3.816 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.888 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.888 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.376 0.108 0.792 0.18 ; 
RECT 0.72 0.504 1.176 0.576 ; 
RECT 0.72 0.108 0.792 0.972 ; 
RECT 0.376 0.9 0.792 0.972 ; 
END 
END BUFx12_ASAP7_75t_R 

MACRO BUFx12f_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN BUFx12f_ASAP7_75t_R 0 0 ; 
SIZE 0.648 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.24 0.108 3.816 0.18 ; 
RECT 3.744 0.108 3.816 0.972 ; 
RECT 1.24 0.9 3.816 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.888 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.888 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.376 0.108 1.116 0.18 ; 
RECT 1.044 0.504 1.244 0.576 ; 
RECT 1.044 0.108 1.116 0.972 ; 
RECT 0.376 0.9 1.116 0.972 ; 
END 
END BUFx12f_ASAP7_75t_R 

MACRO BUFx4_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN BUFx4_ASAP7_75t_R 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.124 0.288 0.292 0.36 ; 
RECT 0.22 0.288 0.292 0.792 ; 
RECT 0.128 0.72 0.292 0.792 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.58 0.144 1.428 0.216 ; 
RECT 1.356 0.144 1.428 0.936 ; 
RECT 0.58 0.864 1.428 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.148 0.108 0.456 0.18 ; 
RECT 0.384 0.504 1.256 0.576 ; 
RECT 0.384 0.108 0.456 0.972 ; 
RECT 0.148 0.9 0.456 0.972 ; 
END 
END BUFx4_ASAP7_75t_R 

MACRO BUFx6f_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN BUFx6f_ASAP7_75t_R 0 0 ; 
SIZE 2.592 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.268 0.36 0.812 ; 
RECT 0.176 0.74 0.36 0.812 ; 
RECT 0.288 0.268 0.48 0.34 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.024 0.108 2.524 0.18 ; 
RECT 2.444 0.108 2.524 0.972 ; 
RECT 1.024 0.9 2.524 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.592 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.592 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.108 0.796 0.18 ; 
RECT 0.716 0.516 1.244 0.588 ; 
RECT 0.716 0.108 0.796 0.972 ; 
RECT 0.16 0.9 0.796 0.972 ; 
END 
END BUFx6f_ASAP7_75t_R 

MACRO BUFx8_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN BUFx8_ASAP7_75t_R 0 0 ; 
SIZE 3.024 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.288 0.36 0.792 ; 
RECT 0.164 0.72 0.36 0.792 ; 
RECT 0.288 0.288 0.5 0.36 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.024 0.144 2.954 0.216 ; 
RECT 2.882 0.144 2.954 0.936 ; 
RECT 1.024 0.864 2.954 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.024 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.024 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.108 0.79 0.18 ; 
RECT 0.718 0.508 1.244 0.58 ; 
RECT 0.718 0.108 0.79 0.972 ; 
RECT 0.16 0.9 0.79 0.972 ; 
END 
END BUFx8_ASAP7_75t_R 

MACRO DECAPx1_ASAP7_75t 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DECAPx1_ASAP7_75t 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.864 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.864 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.292 0.348 0.488 0.42 ; 
RECT 0.292 0.348 0.364 0.6 ; 
RECT 0.564 0.484 0.636 0.772 ; 
RECT 0.376 0.7 0.636 0.772 ; 
RECT 0.992 1.044 1.296 1.116 ; 
RECT 0.992 -0.009 1.296 0.036 ; 
END 
END DECAPx1_ASAP7_75t 

MACRO DECAPxp33_ASAP7_75t 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DECAPxp33_ASAP7_75t 0 0 ; 
SIZE 0.648 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.648 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.648 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.088 0.108 0.272 0.18 ; 
RECT 0.088 0.108 0.16 0.788 ; 
RECT 0.088 0.716 0.312 0.788 ; 
RECT 0.336 0.292 0.56 0.364 ; 
RECT 0.488 0.292 0.56 0.972 ; 
RECT 0.376 0.9 0.56 0.972 ; 
END 
END DECAPxp33_ASAP7_75t 

MACRO DFFHQNx1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DFFHQNx1_ASAP7_75t_R 0 0 ; 
SIZE 4.32 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 4.048 0.108 4.252 0.18 ; 
RECT 4.18 0.108 4.252 0.972 ; 
RECT 4.048 0.9 4.252 0.972 ; 
END 
END QN 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.32 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.32 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.664 0.404 2.736 0.668 ; 
RECT 2.536 0.108 2.952 0.18 ; 
RECT 3.312 0.468 3.384 0.692 ; 
RECT 2.88 0.62 3.384 0.692 ; 
RECT 2.88 0.108 2.952 0.968 ; 
RECT 2.752 0.896 2.952 0.968 ; 
RECT 3.096 0.108 3.6 0.18 ; 
RECT 3.096 0.108 3.168 0.476 ; 
RECT 3.528 0.108 3.6 0.968 ; 
RECT 3.4 0.896 3.6 0.968 ; 
RECT 3.96 0.36 4.032 0.668 ; 
LAYER M2 ; 
RECT 0.704 0.72 2.108 0.792 ; 
RECT 0.076 0.576 2.736 0.648 ; 
RECT 2.88 0.576 4.052 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.96 0.576 4.032 0.648 ; 
END 
END DFFHQNx1_ASAP7_75t_R 

MACRO DFFHQNx2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DFFHQNx2_ASAP7_75t_R 0 0 ; 
SIZE 4.536 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 4.048 0.144 4.468 0.216 ; 
RECT 4.396 0.144 4.468 0.936 ; 
RECT 4.048 0.864 4.468 0.936 ; 
END 
END QN 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.536 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.536 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.664 0.404 2.736 0.668 ; 
RECT 2.536 0.108 2.952 0.18 ; 
RECT 3.312 0.468 3.384 0.692 ; 
RECT 2.88 0.62 3.384 0.692 ; 
RECT 2.88 0.108 2.952 0.968 ; 
RECT 2.752 0.896 2.952 0.968 ; 
RECT 3.096 0.108 3.6 0.18 ; 
RECT 3.096 0.108 3.168 0.476 ; 
RECT 3.528 0.108 3.6 0.968 ; 
RECT 3.4 0.896 3.6 0.968 ; 
RECT 3.96 0.36 4.032 0.668 ; 
LAYER M2 ; 
RECT 0.704 0.72 2.108 0.792 ; 
RECT 0.076 0.576 2.736 0.648 ; 
RECT 2.88 0.576 4.052 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.96 0.576 4.032 0.648 ; 
END 
END DFFHQNx2_ASAP7_75t_R 

MACRO DFFHQNx3_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DFFHQNx3_ASAP7_75t_R 0 0 ; 
SIZE 4.752 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 4.052 0.144 4.684 0.216 ; 
RECT 4.612 0.144 4.684 0.936 ; 
RECT 4.052 0.864 4.684 0.936 ; 
END 
END QN 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.752 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.752 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.664 0.404 2.736 0.668 ; 
RECT 2.536 0.108 2.952 0.18 ; 
RECT 3.312 0.468 3.384 0.692 ; 
RECT 2.88 0.62 3.384 0.692 ; 
RECT 2.88 0.108 2.952 0.968 ; 
RECT 2.752 0.896 2.952 0.968 ; 
RECT 3.096 0.108 3.6 0.18 ; 
RECT 3.096 0.108 3.168 0.476 ; 
RECT 3.528 0.108 3.6 0.968 ; 
RECT 3.4 0.896 3.6 0.968 ; 
RECT 3.96 0.496 4.032 0.668 ; 
LAYER M2 ; 
RECT 0.704 0.72 2.108 0.792 ; 
RECT 0.076 0.576 2.736 0.648 ; 
RECT 2.88 0.576 4.052 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.96 0.576 4.032 0.648 ; 
END 
END DFFHQNx3_ASAP7_75t_R 

MACRO DFFHQNx4_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DFFHQNx4_ASAP7_75t_R 0 0 ; 
SIZE 6.48 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.268 0.332 0.812 ; 
RECT 0.26 0.74 0.48 0.812 ; 
RECT 0.26 0.268 0.492 0.34 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 5.56 0.108 6.412 0.18 ; 
RECT 6.332 0.108 6.412 0.972 ; 
RECT 5.56 0.9 6.412 0.972 ; 
END 
END QN 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 6.48 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 6.48 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.388 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.376 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.664 0.404 2.736 0.668 ; 
RECT 2.536 0.108 2.952 0.18 ; 
RECT 3.312 0.468 3.384 0.692 ; 
RECT 2.88 0.62 3.384 0.692 ; 
RECT 2.88 0.108 2.952 0.968 ; 
RECT 2.752 0.896 2.952 0.968 ; 
RECT 3.096 0.108 3.6 0.18 ; 
RECT 3.096 0.108 3.168 0.476 ; 
RECT 3.528 0.108 3.6 0.968 ; 
RECT 3.4 0.896 3.6 0.968 ; 
RECT 3.96 0.488 4.032 0.668 ; 
RECT 4.048 0.152 4.236 0.224 ; 
RECT 4.164 0.508 4.916 0.58 ; 
RECT 4.164 0.152 4.236 0.936 ; 
RECT 4.048 0.864 4.236 0.936 ; 
RECT 4.48 0.152 5.112 0.224 ; 
RECT 5.04 0.508 6.212 0.58 ; 
RECT 5.04 0.152 5.112 0.936 ; 
RECT 4.696 0.864 5.112 0.936 ; 
LAYER M2 ; 
RECT 0.724 0.72 2.088 0.792 ; 
RECT 0.076 0.576 2.736 0.648 ; 
RECT 2.88 0.576 4.032 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.312 0.576 3.384 0.648 ; 
RECT 3.96 0.576 4.032 0.648 ; 
END 
END DFFHQNx4_ASAP7_75t_R 

MACRO DFFLQNx1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DFFLQNx1_ASAP7_75t_R 0 0 ; 
SIZE 4.32 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 4.048 0.108 4.252 0.18 ; 
RECT 4.18 0.108 4.252 0.972 ; 
RECT 4.048 0.9 4.252 0.972 ; 
END 
END QN 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.32 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.32 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.5 0.508 0.812 0.58 ; 
RECT 0.74 0.508 0.812 0.792 ; 
RECT 0.58 0.72 0.812 0.792 ; 
RECT 0.592 0.108 0.956 0.18 ; 
RECT 0.884 0.108 0.956 0.972 ; 
RECT 0.592 0.9 0.956 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.664 0.404 2.736 0.668 ; 
RECT 2.536 0.108 2.952 0.18 ; 
RECT 3.312 0.468 3.384 0.692 ; 
RECT 2.88 0.62 3.384 0.692 ; 
RECT 2.88 0.108 2.952 0.968 ; 
RECT 2.752 0.896 2.952 0.968 ; 
RECT 3.096 0.108 3.6 0.18 ; 
RECT 3.096 0.108 3.168 0.476 ; 
RECT 3.528 0.108 3.6 0.968 ; 
RECT 3.4 0.896 3.6 0.968 ; 
RECT 3.96 0.36 4.032 0.668 ; 
LAYER M2 ; 
RECT 0.076 0.72 2.108 0.792 ; 
RECT 0.864 0.576 2.736 0.648 ; 
RECT 2.88 0.576 4.052 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.72 0.148 0.792 ; 
RECT 0.6 0.72 0.672 0.792 ; 
RECT 0.884 0.576 0.956 0.648 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.96 0.576 4.032 0.648 ; 
END 
END DFFLQNx1_ASAP7_75t_R 

MACRO DFFLQNx2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DFFLQNx2_ASAP7_75t_R 0 0 ; 
SIZE 4.536 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.296 0.268 0.368 0.8 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.144 1.16 0.8 ; 
RECT 1.088 0.144 1.272 0.216 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 4.048 0.144 4.46 0.216 ; 
RECT 4.388 0.144 4.46 0.936 ; 
RECT 4.052 0.864 4.46 0.936 ; 
END 
END QN 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.536 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.536 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.504 0.476 0.576 0.812 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.664 0.404 2.736 0.668 ; 
RECT 2.536 0.108 2.952 0.18 ; 
RECT 3.312 0.468 3.384 0.692 ; 
RECT 2.88 0.62 3.384 0.692 ; 
RECT 2.88 0.108 2.952 0.968 ; 
RECT 2.752 0.896 2.952 0.968 ; 
RECT 3.096 0.108 3.6 0.18 ; 
RECT 3.096 0.108 3.168 0.476 ; 
RECT 3.528 0.108 3.6 0.968 ; 
RECT 3.4 0.896 3.6 0.968 ; 
RECT 3.96 0.36 4.032 0.668 ; 
LAYER M2 ; 
RECT 0.056 0.72 2.108 0.792 ; 
RECT 0.716 0.576 2.736 0.648 ; 
RECT 2.88 0.576 4.052 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.72 0.148 0.792 ; 
RECT 0.504 0.72 0.576 0.792 ; 
RECT 0.724 0.576 0.796 0.648 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.96 0.576 4.032 0.648 ; 
END 
END DFFLQNx2_ASAP7_75t_R 

MACRO DFFLQNx3_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DFFLQNx3_ASAP7_75t_R 0 0 ; 
SIZE 4.752 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.412 0.576 0.792 ; 
RECT 0.404 0.72 0.576 0.792 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 4.044 0.144 4.684 0.216 ; 
RECT 4.612 0.144 4.684 0.936 ; 
RECT 4.048 0.864 4.684 0.936 ; 
END 
END QN 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.752 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.752 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.26 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.392 0.108 0.796 0.18 ; 
RECT 0.392 0.108 0.464 0.332 ; 
RECT 0.3 0.26 0.464 0.332 ; 
RECT 0.3 0.26 0.372 0.488 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.664 0.404 2.736 0.668 ; 
RECT 2.536 0.108 2.952 0.18 ; 
RECT 3.312 0.468 3.384 0.692 ; 
RECT 2.88 0.62 3.384 0.692 ; 
RECT 2.88 0.108 2.952 0.968 ; 
RECT 2.752 0.896 2.952 0.968 ; 
RECT 3.096 0.108 3.6 0.18 ; 
RECT 3.096 0.108 3.168 0.476 ; 
RECT 3.528 0.108 3.6 0.968 ; 
RECT 3.4 0.896 3.6 0.968 ; 
RECT 3.96 0.36 4.032 0.668 ; 
RECT 4.176 0.36 4.248 0.668 ; 
RECT 4.392 0.36 4.464 0.668 ; 
LAYER M2 ; 
RECT 0.708 0.72 2.108 0.792 ; 
RECT 0.076 0.576 2.736 0.648 ; 
RECT 2.88 0.576 4.484 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.96 0.576 4.032 0.648 ; 
RECT 4.176 0.576 4.248 0.648 ; 
RECT 4.392 0.576 4.464 0.648 ; 
END 
END DFFLQNx3_ASAP7_75t_R 

MACRO DFFLQNx4_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DFFLQNx4_ASAP7_75t_R 0 0 ; 
SIZE 4.968 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.288 0.332 0.684 ; 
RECT 0.26 0.288 0.452 0.36 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.144 1.16 0.812 ; 
RECT 1.088 0.144 1.272 0.216 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 3.812 0.144 4.9 0.216 ; 
RECT 4.828 0.144 4.9 0.936 ; 
RECT 3.812 0.864 4.9 0.936 ; 
END 
END QN 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.968 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.968 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.452 0.584 0.524 0.812 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.664 0.404 2.736 0.668 ; 
RECT 2.536 0.108 2.952 0.18 ; 
RECT 3.312 0.468 3.384 0.692 ; 
RECT 2.88 0.62 3.384 0.692 ; 
RECT 2.88 0.108 2.952 0.968 ; 
RECT 2.752 0.896 2.952 0.968 ; 
RECT 3.096 0.108 3.6 0.18 ; 
RECT 3.096 0.108 3.168 0.476 ; 
RECT 3.528 0.108 3.6 0.968 ; 
RECT 3.4 0.896 3.6 0.968 ; 
RECT 3.96 0.36 4.032 0.668 ; 
LAYER M2 ; 
RECT 0.076 0.72 2.108 0.792 ; 
RECT 0.724 0.576 2.736 0.648 ; 
RECT 2.88 0.576 4.048 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.72 0.148 0.792 ; 
RECT 0.452 0.72 0.524 0.792 ; 
RECT 0.724 0.576 0.796 0.648 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.96 0.576 4.032 0.648 ; 
END 
END DFFLQNx4_ASAP7_75t_R 

MACRO DHLx1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DHLx1_ASAP7_75t_R 0 0 ; 
SIZE 3.24 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN Q 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.968 0.108 3.168 0.18 ; 
RECT 3.096 0.108 3.168 0.972 ; 
RECT 2.968 0.9 3.168 0.972 ; 
END 
END Q 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.24 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.24 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.544 0.508 0.788 0.58 ; 
RECT 0.716 0.508 0.788 0.792 ; 
RECT 0.58 0.72 0.788 0.792 ; 
RECT 0.592 0.108 0.932 0.18 ; 
RECT 0.86 0.108 0.932 0.972 ; 
RECT 0.592 0.9 0.932 0.972 ; 
RECT 1.26 0.5 1.468 0.572 ; 
RECT 1.26 0.5 1.332 0.812 ; 
RECT 1.608 0.48 1.68 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.656 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.32 0.56 ; 
RECT 1.8 0.108 1.872 0.84 ; 
RECT 1.444 0.768 1.872 0.84 ; 
RECT 2.016 0.108 2.52 0.18 ; 
RECT 2.016 0.108 2.088 0.388 ; 
RECT 2.448 0.108 2.52 0.972 ; 
RECT 2.32 0.9 2.52 0.972 ; 
RECT 2.732 0.268 2.804 0.58 ; 
RECT 2.732 0.508 2.972 0.58 ; 
LAYER M2 ; 
RECT 0.84 0.576 1.7 0.648 ; 
RECT 0.076 0.72 2.172 0.792 ; 
RECT 1.776 0.288 3.004 0.36 ; 
LAYER V1 ; 
RECT 0.076 0.72 0.148 0.792 ; 
RECT 0.6 0.72 0.672 0.792 ; 
RECT 0.86 0.576 0.932 0.648 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.608 0.576 1.68 0.648 ; 
RECT 1.8 0.288 1.872 0.36 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.732 0.288 2.804 0.36 ; 
END 
END DHLx1_ASAP7_75t_R 

MACRO DHLx2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DHLx2_ASAP7_75t_R 0 0 ; 
SIZE 3.456 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.256 0.288 0.328 0.668 ; 
RECT 0.416 0.14 0.488 0.36 ; 
RECT 0.256 0.288 0.488 0.36 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.824 ; 
END 
END D 
PIN Q 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.972 0.144 3.4 0.216 ; 
RECT 3.328 0.144 3.4 0.936 ; 
RECT 2.964 0.864 3.4 0.936 ; 
END 
END Q 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.456 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.456 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.476 0.64 0.792 ; 
RECT 0.432 0.72 0.64 0.792 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 2.88 0.36 2.952 0.668 ; 
RECT 3.096 0.36 3.168 0.668 ; 
LAYER M2 ; 
RECT 0.708 0.576 1.668 0.648 ; 
RECT 0.064 0.72 2.104 0.792 ; 
RECT 1.792 0.576 3.192 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.72 0.148 0.792 ; 
RECT 0.496 0.72 0.568 0.792 ; 
RECT 0.724 0.576 0.796 0.648 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 1.8 0.576 1.872 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.88 0.576 2.952 0.648 ; 
RECT 3.096 0.576 3.168 0.648 ; 
END 
END DHLx2_ASAP7_75t_R 

MACRO DHLx3_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DHLx3_ASAP7_75t_R 0 0 ; 
SIZE 3.888 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.288 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.36 ; 
RECT 0.26 0.288 0.492 0.36 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.144 0.276 1.216 0.812 ; 
END 
END D 
PIN Q 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.968 0.108 3.816 0.18 ; 
RECT 3.744 0.108 3.816 0.972 ; 
RECT 2.968 0.9 3.816 0.972 ; 
END 
END Q 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.888 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.888 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.552 0.488 0.624 0.668 ; 
RECT 0.596 0.108 0.8 0.18 ; 
RECT 0.728 0.108 0.8 0.972 ; 
RECT 0.596 0.9 0.8 0.972 ; 
RECT 1.368 0.432 1.44 0.668 ; 
RECT 1.74 0.544 1.912 0.616 ; 
RECT 1.74 0.544 1.812 0.812 ; 
RECT 1.556 0.36 2.088 0.432 ; 
RECT 2.012 0.36 2.088 0.804 ; 
RECT 2.012 0.732 2.452 0.804 ; 
RECT 2.264 0.66 2.336 0.876 ; 
RECT 1.556 0.36 1.628 0.908 ; 
RECT 1.472 0.836 1.628 0.908 ; 
RECT 2.228 0.36 2.628 0.432 ; 
RECT 2.556 0.136 2.628 0.94 ; 
RECT 2.756 0.492 3.156 0.564 ; 
RECT 2.756 0.492 2.828 0.812 ; 
LAYER M2 ; 
RECT 0.072 0.576 1.664 0.648 ; 
RECT 0.708 0.72 1.896 0.792 ; 
RECT 2.264 0.72 2.848 0.792 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.552 0.576 0.624 0.648 ; 
RECT 0.728 0.72 0.8 0.792 ; 
RECT 1.368 0.576 1.44 0.648 ; 
RECT 1.74 0.72 1.812 0.792 ; 
RECT 2.264 0.72 2.336 0.792 ; 
RECT 2.756 0.72 2.828 0.792 ; 
END 
END DHLx3_ASAP7_75t_R 

MACRO DLLx1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DLLx1_ASAP7_75t_R 0 0 ; 
SIZE 3.24 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN Q 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.94 0.108 3.168 0.18 ; 
RECT 3.096 0.108 3.168 0.972 ; 
RECT 2.968 0.9 3.168 0.972 ; 
END 
END Q 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.24 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.24 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.572 0.488 0.644 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.264 0.5 1.468 0.572 ; 
RECT 1.264 0.5 1.336 0.812 ; 
RECT 1.608 0.48 1.68 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.656 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.32 0.56 ; 
RECT 1.8 0.108 1.872 0.84 ; 
RECT 1.444 0.768 1.872 0.84 ; 
RECT 2.016 0.108 2.52 0.18 ; 
RECT 2.016 0.108 2.088 0.388 ; 
RECT 2.448 0.108 2.52 0.972 ; 
RECT 2.32 0.9 2.52 0.972 ; 
RECT 2.712 0.268 2.784 0.58 ; 
RECT 2.712 0.508 2.972 0.58 ; 
LAYER M2 ; 
RECT 0.076 0.576 1.7 0.648 ; 
RECT 0.682 0.72 2.172 0.792 ; 
RECT 1.776 0.288 3.004 0.36 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.572 0.576 0.644 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.264 0.72 1.336 0.792 ; 
RECT 1.608 0.576 1.68 0.648 ; 
RECT 1.8 0.288 1.872 0.36 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.712 0.288 2.784 0.36 ; 
END 
END DLLx1_ASAP7_75t_R 

MACRO DLLx2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DLLx2_ASAP7_75t_R 0 0 ; 
SIZE 3.456 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.412 0.332 0.792 ; 
RECT 0.26 0.72 0.424 0.792 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN Q 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.752 0.108 3.388 0.18 ; 
RECT 3.316 0.108 3.388 0.972 ; 
RECT 2.752 0.9 3.388 0.972 ; 
END 
END Q 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.456 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.456 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.392 0.64 0.696 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.544 0.416 ; 
RECT 2.472 0.344 2.544 0.968 ; 
RECT 2.304 0.896 2.544 0.968 ; 
RECT 3.096 0.36 3.168 0.668 ; 
LAYER M2 ; 
RECT 0.076 0.576 1.656 0.648 ; 
RECT 0.724 0.72 2.108 0.792 ; 
RECT 1.8 0.576 3.2 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 1.8 0.576 1.872 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 3.096 0.576 3.168 0.648 ; 
END 
END DLLx2_ASAP7_75t_R 

MACRO DLLx3_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN DLLx3_ASAP7_75t_R 0 0 ; 
SIZE 3.672 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.088 0.268 1.16 0.812 ; 
END 
END D 
PIN Q 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.968 0.144 3.604 0.216 ; 
RECT 3.528 0.144 3.604 0.936 ; 
RECT 2.968 0.864 3.604 0.936 ; 
END 
END Q 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.672 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.672 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.26 0.492 1.468 0.564 ; 
RECT 1.26 0.492 1.332 0.812 ; 
RECT 1.584 0.432 1.656 0.668 ; 
RECT 2.016 0.66 2.088 0.812 ; 
RECT 1.672 0.108 1.872 0.18 ; 
RECT 1.8 0.488 2.312 0.56 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.456 0.9 1.872 0.972 ; 
RECT 2.34 0.18 2.412 0.416 ; 
RECT 1.984 0.344 2.524 0.416 ; 
RECT 2.444 0.344 2.524 0.968 ; 
RECT 2.304 0.896 2.524 0.968 ; 
RECT 2.66 0.508 3.416 0.58 ; 
RECT 2.66 0.508 2.74 0.796 ; 
LAYER M2 ; 
RECT 0.076 0.576 1.672 0.648 ; 
RECT 0.704 0.72 2.108 0.792 ; 
RECT 1.8 0.576 2.792 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.26 0.72 1.332 0.792 ; 
RECT 1.584 0.576 1.656 0.648 ; 
RECT 1.8 0.576 1.872 0.648 ; 
RECT 2.016 0.72 2.088 0.792 ; 
RECT 2.664 0.576 2.736 0.648 ; 
END 
END DLLx3_ASAP7_75t_R 

MACRO FILLER_ASAP7_75t 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN FILLER_ASAP7_75t 0 0 ; 
SIZE 0.432 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.432 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.432 0.036 ; 
END 
END vss! 
END FILLER_ASAP7_75t 
####################################
MACRO FILLER_TEST_ASAP7_75t
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN FILLER_TEST_ASAP7_75t 0 0 ; 
SIZE 0.432 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.432 1.116 ;
END
END vdd!

PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.432 0.036 ; 
END
END vss!
END FILLER_TEST_ASAP7_75t 

MACRO FILLER_TEST1_ASAP7_75t
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN FILLER_TEST1_ASAP7_75t 0 0 ; 
SIZE 0.216 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.216 1.116 ;
END
END vdd!

PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.216 0.036 ; 
END
END vss!
END FILLER_TEST1_ASAP7_75t 
####################################
MACRO HB1xp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN HB1xp67_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.024 0.144 1.224 0.216 ; 
RECT 1.152 0.144 1.224 0.972 ; 
RECT 1.024 0.9 1.224 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.376 0.108 0.576 0.18 ; 
RECT 0.504 0.504 0.96 0.576 ; 
RECT 0.504 0.108 0.576 0.972 ; 
RECT 0.376 0.9 0.576 0.972 ; 
END 
END HB1xp67_ASAP7_75t_R 

MACRO HB2xp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN HB2xp67_ASAP7_75t_R 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.224 0.256 0.296 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.24 0.144 1.44 0.216 ; 
RECT 1.368 0.144 1.44 0.936 ; 
RECT 1.24 0.864 1.44 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.592 0.108 0.792 0.18 ; 
RECT 0.72 0.504 1.232 0.576 ; 
RECT 0.72 0.108 0.792 0.972 ; 
RECT 0.592 0.9 0.792 0.972 ; 
END 
END HB2xp67_ASAP7_75t_R 

MACRO HB3xp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN HB3xp67_ASAP7_75t_R 0 0 ; 
SIZE 1.728 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.456 0.144 1.656 0.216 ; 
RECT 1.584 0.144 1.656 0.936 ; 
RECT 1.456 0.864 1.656 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.728 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.728 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.808 0.108 1.008 0.18 ; 
RECT 0.936 0.468 1.44 0.54 ; 
RECT 0.936 0.108 1.008 0.972 ; 
RECT 0.808 0.9 1.008 0.972 ; 
END 
END HB3xp67_ASAP7_75t_R 

MACRO HB4xp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN HB4xp67_ASAP7_75t_R 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.224 0.288 0.296 0.792 ; 
RECT 0.14 0.72 0.296 0.792 ; 
RECT 0.224 0.288 0.476 0.36 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.24 0.144 1.44 0.216 ; 
RECT 1.368 0.144 1.44 0.936 ; 
RECT 1.24 0.864 1.44 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.108 0.752 0.18 ; 
RECT 0.68 0.404 1.2 0.476 ; 
RECT 0.68 0.108 0.752 0.972 ; 
RECT 0.16 0.9 0.752 0.972 ; 
END 
END HB4xp67_ASAP7_75t_R 

MACRO ICGNx1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN -0.054 0 ; 
FOREIGN ICGNx1_ASAP7_75t_R 0.216 0 ; 
SIZE 4.104 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.268 0.268 0.34 0.72 ; 
RECT 0.268 0.268 0.58 0.34 ; 
END 
END CLK 
PIN EN 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.368 0.268 1.44 0.972 ; 
RECT 1.26 0.9 1.44 0.972 ; 
RECT 1.368 0.268 1.564 0.34 ; 
END 
END EN 
PIN GCLKN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 3.612 0.108 4.248 0.18 ; 
RECT 4.176 0.108 4.248 0.972 ; 
RECT 3.392 0.9 4.248 0.972 ; 
END 
END GCLKN 
PIN SE 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.956 0.268 1.16 0.34 ; 
RECT 1.088 0.268 1.16 0.972 ; 
RECT 0.924 0.9 1.16 0.972 ; 
END 
END SE 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.32 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.32 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.26 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.452 0.584 0.524 0.812 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.004 0.108 1.592 0.18 ; 
RECT 1.584 0.46 1.656 0.812 ; 
RECT 1.8 0.432 1.872 0.668 ; 
RECT 2.232 0.66 2.304 0.812 ; 
RECT 1.888 0.108 2.088 0.18 ; 
RECT 2.016 0.488 2.528 0.56 ; 
RECT 2.016 0.108 2.088 0.972 ; 
RECT 1.672 0.9 2.088 0.972 ; 
RECT 2.556 0.18 2.628 0.416 ; 
RECT 2.2 0.344 2.76 0.416 ; 
RECT 2.688 0.496 3.192 0.568 ; 
RECT 2.688 0.344 2.76 0.968 ; 
RECT 2.52 0.896 2.76 0.968 ; 
RECT 2.932 0.304 3.972 0.376 ; 
RECT 3.528 0.476 3.6 0.72 ; 
RECT 3.96 0.476 4.032 0.72 ; 
RECT 3.256 0.648 4.032 0.72 ; 
RECT 3.256 0.648 3.328 0.82 ; 
LAYER M2 ; 
RECT 0.724 0.576 1.968 0.648 ; 
RECT 0.076 0.72 3.388 0.792 ; 
LAYER V1 ; 
RECT 0.076 0.72 0.148 0.792 ; 
RECT 0.452 0.72 0.524 0.792 ; 
RECT 0.724 0.576 0.796 0.648 ; 
RECT 1.584 0.72 1.656 0.792 ; 
RECT 1.8 0.576 1.872 0.648 ; 
RECT 2.232 0.72 2.304 0.792 ; 
RECT 3.256 0.72 3.328 0.792 ; 
END 
END ICGNx1_ASAP7_75t_R 

MACRO ICGNx2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN ICGNx2_ASAP7_75t_R 0 0 ; 
SIZE 5.4 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN EN 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.332 0.252 1.404 0.936 ; 
RECT 1.332 0.864 1.496 0.936 ; 
RECT 1.332 0.252 1.504 0.324 ; 
END 
END EN 
PIN GCLKN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 4.824 0.108 4.896 0.972 ; 
RECT 4.696 0.108 5.024 0.18 ; 
RECT 4.696 0.9 5.024 0.972 ; 
END 
END GCLKN 
PIN SE 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.984 0.252 1.16 0.324 ; 
RECT 1.088 0.252 1.16 0.936 ; 
RECT 0.896 0.864 1.16 0.936 ; 
END 
END SE 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 5.4 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 5.4 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.024 0.108 1.568 0.18 ; 
RECT 1.476 0.492 1.684 0.564 ; 
RECT 1.476 0.492 1.548 0.672 ; 
RECT 1.8 0.432 1.872 0.792 ; 
RECT 1.668 0.72 1.872 0.792 ; 
RECT 2.232 0.66 2.304 0.812 ; 
RECT 2.448 0.484 2.52 0.668 ; 
RECT 1.888 0.108 2.088 0.18 ; 
RECT 2.32 0.108 2.736 0.18 ; 
RECT 2.016 0.312 2.736 0.384 ; 
RECT 3.096 0.468 3.168 0.692 ; 
RECT 2.664 0.62 3.168 0.692 ; 
RECT 2.016 0.108 2.088 0.936 ; 
RECT 1.672 0.864 2.088 0.936 ; 
RECT 2.664 0.108 2.736 0.968 ; 
RECT 2.536 0.896 2.736 0.968 ; 
RECT 2.88 0.108 3.384 0.18 ; 
RECT 2.88 0.108 2.952 0.476 ; 
RECT 3.312 0.108 3.384 0.968 ; 
RECT 3.184 0.896 3.384 0.968 ; 
RECT 3.636 0.136 3.708 0.38 ; 
RECT 3.676 0.556 3.748 0.812 ; 
RECT 3.892 0.288 3.964 0.812 ; 
RECT 4.048 0.108 4.248 0.18 ; 
RECT 4.176 0.272 4.68 0.344 ; 
RECT 4.608 0.272 4.68 0.812 ; 
RECT 4.176 0.108 4.248 0.972 ; 
RECT 4.048 0.9 4.248 0.972 ; 
RECT 5.04 0.268 5.112 0.812 ; 
LAYER M2 ; 
RECT 0.076 0.576 2.52 0.648 ; 
RECT 2.664 0.576 3.748 0.648 ; 
RECT 0.704 0.72 3.984 0.792 ; 
RECT 3.616 0.288 4.268 0.36 ; 
RECT 4.58 0.576 5.128 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 1.476 0.576 1.548 0.648 ; 
RECT 1.688 0.72 1.76 0.792 ; 
RECT 2.232 0.72 2.304 0.792 ; 
RECT 2.448 0.576 2.52 0.648 ; 
RECT 2.664 0.576 2.736 0.648 ; 
RECT 3.636 0.288 3.708 0.36 ; 
RECT 3.676 0.576 3.748 0.648 ; 
RECT 3.892 0.72 3.964 0.792 ; 
RECT 4.176 0.288 4.248 0.36 ; 
RECT 4.608 0.576 4.68 0.648 ; 
RECT 5.04 0.576 5.112 0.648 ; 
END 
END ICGNx2_ASAP7_75t_R 

MACRO ICGx2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN ICGx2_ASAP7_75t_R 0 0 ; 
SIZE 5.832 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.28 0.332 0.8 ; 
RECT 0.26 0.728 0.48 0.8 ; 
RECT 0.408 0.728 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.352 ; 
RECT 0.26 0.28 0.492 0.352 ; 
END 
END CLK 
PIN EN 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.932 0.144 1.108 0.216 ; 
RECT 1.036 0.144 1.108 0.352 ; 
RECT 1.036 0.28 1.224 0.352 ; 
RECT 1.152 0.28 1.224 0.648 ; 
END 
END EN 
PIN GCLK 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 5.128 0.144 5.764 0.216 ; 
RECT 5.692 0.144 5.764 0.936 ; 
RECT 5.128 0.864 5.764 0.936 ; 
END 
END GCLK 
PIN SE 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.356 0.284 1.428 0.616 ; 
END 
END SE 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 5.832 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 5.832 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.24 0.108 1.572 0.18 ; 
RECT 1.5 0.436 1.672 0.508 ; 
RECT 1.5 0.108 1.572 0.828 ; 
RECT 1.024 0.756 1.572 0.828 ; 
RECT 1.672 0.108 1.876 0.18 ; 
RECT 1.804 0.504 2.24 0.576 ; 
RECT 1.804 0.108 1.876 0.972 ; 
RECT 1.672 0.9 1.876 0.972 ; 
RECT 2.34 0.492 2.548 0.564 ; 
RECT 2.34 0.492 2.412 0.668 ; 
RECT 2.664 0.472 2.736 0.792 ; 
RECT 2.532 0.72 2.736 0.792 ; 
RECT 3.744 0.528 3.816 0.688 ; 
RECT 2.752 0.108 3.948 0.18 ; 
RECT 2.88 0.488 3.404 0.56 ; 
RECT 2.88 0.108 2.952 0.972 ; 
RECT 2.536 0.9 2.952 0.972 ; 
RECT 3.064 0.344 4.036 0.416 ; 
RECT 3.552 0.344 3.624 0.968 ; 
RECT 3.384 0.896 3.624 0.968 ; 
RECT 4.316 0.632 4.388 0.812 ; 
RECT 4.688 0.108 4.864 0.18 ; 
RECT 4.792 0.508 5.348 0.58 ; 
RECT 4.792 0.108 4.864 0.972 ; 
RECT 4.48 0.9 4.864 0.972 ; 
LAYER M2 ; 
RECT 0.072 0.576 3.828 0.648 ; 
RECT 0.7 0.72 4.408 0.792 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 2.34 0.576 2.412 0.648 ; 
RECT 2.552 0.72 2.624 0.792 ; 
RECT 3.744 0.576 3.816 0.648 ; 
RECT 4.316 0.72 4.388 0.792 ; 
END 
PROPERTY oaTaper "__DerivedDefaultTaperCG" ; 
END ICGx2_ASAP7_75t_R 

MACRO ICGx3_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN ICGx3_ASAP7_75t_R 0 0 ; 
SIZE 7.344 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.288 0.332 0.936 ; 
RECT 0.26 0.864 0.424 0.936 ; 
RECT 0.42 0.14 0.492 0.36 ; 
RECT 0.26 0.288 0.492 0.36 ; 
END 
END CLK 
PIN EN 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.9 0.576 0.972 0.792 ; 
RECT 0.964 0.136 1.036 0.36 ; 
RECT 0.964 0.288 1.224 0.36 ; 
RECT 1.152 0.288 1.224 0.648 ; 
RECT 0.9 0.576 1.224 0.648 ; 
END 
END EN 
PIN GCLK 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 6.64 0.144 7.272 0.216 ; 
RECT 7.2 0.144 7.272 0.972 ; 
RECT 6.62 0.9 7.272 0.972 ; 
END 
END GCLK 
PIN SE 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.452 0.288 1.656 0.36 ; 
RECT 1.584 0.288 1.656 0.648 ; 
RECT 1.584 0.576 1.752 0.648 ; 
END 
END SE 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 7.344 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 7.344 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.08 0.108 0.276 0.18 ; 
RECT 0.08 0.108 0.152 0.892 ; 
RECT 0.568 0.432 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.024 0.9 2 0.972 ; 
RECT 1.24 0.108 2.092 0.18 ; 
RECT 2.012 0.504 2.972 0.576 ; 
RECT 2.012 0.108 2.092 0.792 ; 
RECT 1.672 0.72 2.092 0.792 ; 
RECT 2.536 0.312 3.168 0.384 ; 
RECT 3.096 0.504 3.56 0.576 ; 
RECT 3.096 0.312 3.168 0.772 ; 
RECT 2.536 0.7 3.168 0.772 ; 
RECT 3.744 0.476 3.816 0.736 ; 
RECT 3.836 0.288 4.032 0.36 ; 
RECT 3.96 0.288 4.032 0.792 ; 
RECT 3.96 0.72 4.104 0.792 ; 
RECT 4.392 0.48 4.464 0.648 ; 
RECT 4.392 0.576 4.596 0.648 ; 
RECT 4.048 0.108 4.276 0.18 ; 
RECT 4.204 0.724 4.7 0.796 ; 
RECT 4.204 0.108 4.276 0.964 ; 
RECT 3.832 0.892 4.276 0.964 ; 
RECT 4.696 0.12 4.896 0.192 ; 
RECT 4.376 0.292 4.896 0.364 ; 
RECT 4.82 0.496 5.348 0.568 ; 
RECT 4.82 0.12 4.896 0.968 ; 
RECT 4.68 0.896 4.896 0.968 ; 
RECT 5.596 0.516 5.78 0.588 ; 
RECT 5.596 0.516 5.668 0.792 ; 
RECT 5.596 0.72 5.884 0.792 ; 
RECT 5.128 0.16 6.104 0.232 ; 
RECT 5.776 0.332 6.192 0.404 ; 
RECT 6.116 0.508 7.076 0.58 ; 
RECT 6.116 0.332 6.192 0.96 ; 
RECT 5.344 0.888 6.192 0.96 ; 
LAYER M2 ; 
RECT 0.08 0.576 4.688 0.648 ; 
RECT 0.724 0.72 5.864 0.792 ; 
LAYER V1 ; 
RECT 0.08 0.576 0.152 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 3.744 0.576 3.816 0.648 ; 
RECT 4.012 0.72 4.084 0.792 ; 
RECT 4.504 0.576 4.576 0.648 ; 
RECT 5.792 0.72 5.864 0.792 ; 
END 
END ICGx3_ASAP7_75t_R 

MACRO INVx11_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx11_ASAP7_75t_R 0 0 ; 
SIZE 2.808 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 2.756 0.18 ; 
RECT 2.684 0.108 2.756 0.972 ; 
RECT 0.376 0.9 2.756 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.808 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.808 0.036 ; 
END 
END vss! 
END INVx11_ASAP7_75t_R 

MACRO INVx13_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx13_ASAP7_75t_R 0 0 ; 
SIZE 3.24 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 3.172 0.18 ; 
RECT 3.1 0.108 3.172 0.972 ; 
RECT 0.376 0.9 3.172 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.24 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.24 0.036 ; 
END 
END vss! 
END INVx13_ASAP7_75t_R 

MACRO INVx1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx1_ASAP7_75t_R 0 0 ; 
SIZE 0.648 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 0.576 0.18 ; 
RECT 0.504 0.108 0.576 0.972 ; 
RECT 0.376 0.9 0.576 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.648 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.648 0.036 ; 
END 
END vss! 
END INVx1_ASAP7_75t_R 

MACRO INVx2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx2_ASAP7_75t_R 0 0 ; 
SIZE 0.864 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 0.788 0.18 ; 
RECT 0.716 0.108 0.788 0.972 ; 
RECT 0.376 0.9 0.788 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.864 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.864 0.036 ; 
END 
END vss! 
END INVx2_ASAP7_75t_R 

MACRO INVx3_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx3_ASAP7_75t_R 0 0 ; 
SIZE 1.08 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 1.004 0.18 ; 
RECT 0.932 0.108 1.004 0.972 ; 
RECT 0.376 0.9 1.004 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.08 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.08 0.036 ; 
END 
END vss! 
END INVx3_ASAP7_75t_R 

MACRO INVx4_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx4_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 1.168 0.18 ; 
RECT 1.096 0.108 1.168 0.972 ; 
RECT 0.376 0.9 1.168 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
END INVx4_ASAP7_75t_R 

MACRO INVx5_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx5_ASAP7_75t_R 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.808 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 1.432 0.18 ; 
RECT 1.36 0.108 1.432 0.972 ; 
RECT 0.376 0.9 1.432 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
END INVx5_ASAP7_75t_R 

MACRO INVx6_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx6_ASAP7_75t_R 0 0 ; 
SIZE 1.728 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.808 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 1.648 0.18 ; 
RECT 1.576 0.108 1.648 0.972 ; 
RECT 0.376 0.9 1.648 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.728 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.728 0.036 ; 
END 
END vss! 
END INVx6_ASAP7_75t_R 

MACRO INVx8_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVx8_ASAP7_75t_R 0 0 ; 
SIZE 2.16 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 2.048 0.18 ; 
RECT 1.976 0.108 2.048 0.972 ; 
RECT 0.376 0.9 2.048 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.16 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.16 0.036 ; 
END 
END vss! 
END INVx8_ASAP7_75t_R 

MACRO INVxp33_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVxp33_ASAP7_75t_R 0 0 ; 
SIZE 0.648 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 0.576 0.18 ; 
RECT 0.504 0.108 0.576 0.972 ; 
RECT 0.376 0.9 0.576 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.648 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.648 0.036 ; 
END 
END vss! 
END INVxp33_ASAP7_75t_R 

MACRO INVxp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN INVxp67_ASAP7_75t_R 0 0 ; 
SIZE 0.648 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 0.576 0.18 ; 
RECT 0.504 0.108 0.576 0.972 ; 
RECT 0.376 0.9 0.576 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.648 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.648 0.036 ; 
END 
END vss! 
END INVxp67_ASAP7_75t_R 

MACRO MAJIxp5_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN MAJIxp5_ASAP7_75t_R 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.22 0.48 1.292 0.648 ; 
RECT 1.112 0.576 1.292 0.648 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.224 0.276 0.296 0.792 ; 
RECT 0.856 0.496 0.928 0.792 ; 
RECT 0.224 0.72 0.928 0.792 ; 
RECT 0.856 0.496 1.008 0.568 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.288 0.576 0.62 ; 
RECT 0.504 0.288 0.72 0.36 ; 
END 
END C 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.028 0.288 1.444 0.36 ; 
RECT 1.372 0.288 1.444 0.792 ; 
RECT 1.028 0.72 1.444 0.792 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.376 0.9 1.352 0.972 ; 
RECT 0.376 0.108 1.352 0.18 ; 
END 
END MAJIxp5_ASAP7_75t_R 

MACRO NAND2x1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NAND2x1_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.244 0.412 0.316 0.812 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.584 0.432 0.9 0.504 ; 
RECT 0.828 0.432 0.9 0.668 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.808 0.252 1.228 0.324 ; 
RECT 1.156 0.252 1.228 0.972 ; 
RECT 0.376 0.9 1.228 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.108 1.136 0.18 ; 
END 
END NAND2x1_ASAP7_75t_R 

MACRO NAND2xp33_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NAND2xp33_ASAP7_75t_R 0 0 ; 
SIZE 0.864 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.412 0.576 0.668 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.572 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.376 0.9 0.796 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.864 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.864 0.036 ; 
END 
END vss! 
END NAND2xp33_ASAP7_75t_R 

MACRO NAND2xp5_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NAND2xp5_ASAP7_75t_R 0 0 ; 
SIZE 0.864 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.136 0.108 0.292 0.18 ; 
RECT 0.22 0.108 0.292 0.812 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.424 0.268 0.576 0.34 ; 
RECT 0.504 0.268 0.576 0.812 ; 
RECT 0.428 0.74 0.576 0.812 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.572 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.376 0.9 0.796 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.864 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.864 0.036 ; 
END 
END vss! 
END NAND2xp5_ASAP7_75t_R 

MACRO NAND2xp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NAND2xp67_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.412 0.36 0.812 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.636 0.432 1.008 0.504 ; 
RECT 0.936 0.432 1.008 0.668 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.808 0.252 1.152 0.324 ; 
RECT 1.08 0.252 1.152 0.972 ; 
RECT 0.592 0.9 1.152 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.108 1.136 0.18 ; 
END 
END NAND2xp67_ASAP7_75t_R 

MACRO NAND3x1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NAND3x1_ASAP7_75t_R 0 0 ; 
SIZE 2.376 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.6 0.432 1.872 0.504 ; 
RECT 1.8 0.432 1.872 0.792 ; 
RECT 1.608 0.72 1.872 0.792 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.984 0.432 1.224 0.504 ; 
RECT 1.152 0.432 1.224 0.792 ; 
RECT 0.972 0.72 1.224 0.792 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.244 0.412 0.316 0.812 ; 
END 
END C 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.672 0.252 2.304 0.324 ; 
RECT 2.232 0.252 2.304 0.972 ; 
RECT 0.808 0.9 2.304 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.376 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.376 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.108 0.704 0.18 ; 
RECT 0.376 0.252 1.352 0.324 ; 
RECT 1.024 0.108 2 0.18 ; 
END 
END NAND3x1_ASAP7_75t_R 

MACRO NAND4xp25_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NAND4xp25_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.288 1.008 0.668 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.268 0.792 0.668 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.268 0.576 0.668 ; 
END 
END C 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.168 0.144 0.36 0.216 ; 
RECT 0.288 0.144 0.36 0.792 ; 
RECT 0.168 0.72 0.36 0.792 ; 
END 
END D 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.024 0.108 1.22 0.18 ; 
RECT 1.148 0.108 1.22 0.936 ; 
RECT 0.16 0.864 1.22 0.936 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
END NAND4xp25_ASAP7_75t_R 

MACRO NAND5xp2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NAND5xp2_ASAP7_75t_R 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.288 0.36 0.8 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.136 0.576 0.8 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.136 0.792 0.8 ; 
END 
END C 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.136 1.008 0.8 ; 
END 
END D 
PIN E 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.152 0.136 1.224 0.8 ; 
END 
END E 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.068 0.108 0.148 0.972 ; 
RECT 0.068 0.108 0.28 0.18 ; 
RECT 0.068 0.9 1.352 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
END NAND5xp2_ASAP7_75t_R 

MACRO NOR2x1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NOR2x1_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.244 0.268 0.316 0.668 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.828 0.412 0.9 0.648 ; 
RECT 0.584 0.576 0.9 0.648 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 1.228 0.18 ; 
RECT 1.156 0.108 1.228 0.828 ; 
RECT 0.808 0.756 1.228 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 1.136 0.972 ; 
END 
END NOR2x1_ASAP7_75t_R 

MACRO NOR2xp33_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NOR2xp33_ASAP7_75t_R 0 0 ; 
SIZE 0.864 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.268 0.292 0.812 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.412 0.576 0.668 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.376 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.572 0.9 0.796 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.864 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.864 0.036 ; 
END 
END vss! 
END NOR2xp33_ASAP7_75t_R 

MACRO NOR2xp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NOR2xp67_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.268 0.36 0.668 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.412 1.008 0.648 ; 
RECT 0.636 0.576 1.008 0.648 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.592 0.108 1.152 0.18 ; 
RECT 1.08 0.108 1.152 0.828 ; 
RECT 0.808 0.756 1.152 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 1.136 0.972 ; 
END 
END NOR2xp67_ASAP7_75t_R 

MACRO NOR3x1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NOR3x1_ASAP7_75t_R 0 0 ; 
SIZE 2.376 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.608 0.288 1.872 0.36 ; 
RECT 1.8 0.288 1.872 0.648 ; 
RECT 1.6 0.576 1.872 0.648 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.972 0.288 1.224 0.36 ; 
RECT 1.152 0.288 1.224 0.648 ; 
RECT 0.984 0.576 1.224 0.648 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.244 0.268 0.316 0.668 ; 
END 
END C 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.808 0.108 2.304 0.18 ; 
RECT 2.232 0.108 2.304 0.828 ; 
RECT 1.672 0.756 2.304 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.376 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.376 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.16 0.9 0.704 0.972 ; 
RECT 0.376 0.756 1.352 0.828 ; 
RECT 1.024 0.9 2 0.972 ; 
END 
END NOR3x1_ASAP7_75t_R 

MACRO NOR4xp25_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NOR4xp25_ASAP7_75t_R 0 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.412 1.008 0.792 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.412 0.792 0.812 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.412 0.576 0.812 ; 
END 
END C 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.168 0.288 0.36 0.36 ; 
RECT 0.288 0.288 0.36 0.936 ; 
RECT 0.168 0.864 0.36 0.936 ; 
END 
END D 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.16 0.144 1.22 0.216 ; 
RECT 1.148 0.144 1.22 0.972 ; 
RECT 1.024 0.9 1.22 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.296 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.296 0.036 ; 
END 
END vss! 
END NOR4xp25_ASAP7_75t_R 

MACRO NOR5xp2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN NOR5xp2_ASAP7_75t_R 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.28 0.36 0.792 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.28 0.576 0.944 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.28 0.792 0.944 ; 
END 
END C 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.28 1.008 0.944 ; 
END 
END D 
PIN E 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.152 0.28 1.224 0.944 ; 
END 
END E 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.068 0.108 0.148 0.972 ; 
RECT 0.068 0.9 0.28 0.972 ; 
RECT 0.068 0.108 1.352 0.18 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
END NOR5xp2_ASAP7_75t_R 

MACRO O2A1Ixp5_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN O2A1Ixp5_ASAP7_75t_R 0 0 ; 
SIZE 1.728 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.232 0.252 0.304 0.812 ; 
RECT 0.232 0.252 1.004 0.324 ; 
RECT 0.932 0.252 1.004 0.684 ; 
RECT 0.796 0.612 1.004 0.684 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.436 0.424 0.508 0.8 ; 
RECT 0.436 0.5 0.64 0.572 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.148 0.392 1.22 0.656 ; 
END 
END B 
PIN C 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.34 0.268 1.508 0.34 ; 
RECT 1.436 0.268 1.508 0.656 ; 
END 
END C 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.256 0.108 1.656 0.18 ; 
RECT 1.58 0.108 1.656 0.972 ; 
RECT 1.456 0.9 1.656 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.728 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.728 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.384 0.9 0.912 0.972 ; 
RECT 0.608 0.108 1.12 0.18 ; 
RECT 0.608 0.756 1.34 0.828 ; 
END 
END O2A1Ixp5_ASAP7_75t_R 

MACRO OA21x2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN OA21x2_ASAP7_75t_R 0 0 ; 
SIZE 1.512 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.116 0.252 0.292 0.324 ; 
RECT 0.22 0.252 0.292 0.972 ; 
RECT 0.12 0.9 0.292 0.972 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.424 0.576 0.812 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.716 0.424 0.788 0.684 ; 
RECT 0.716 0.612 0.956 0.684 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.032 0.108 1.44 0.18 ; 
RECT 1.368 0.108 1.44 0.972 ; 
RECT 1.024 0.9 1.44 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.512 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.512 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.168 0.108 0.696 0.18 ; 
RECT 0.396 0.252 1.224 0.324 ; 
RECT 1.152 0.252 1.224 0.828 ; 
RECT 0.824 0.756 1.224 0.828 ; 
RECT 0.824 0.756 0.896 0.972 ; 
RECT 0.592 0.9 0.896 0.972 ; 
END 
END OA21x2_ASAP7_75t_R 

MACRO OA22x2_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN OA22x2_ASAP7_75t_R 0 0 ; 
SIZE 2.16 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.976 0.412 1.156 0.484 ; 
RECT 1.084 0.412 1.156 0.812 ; 
RECT 0.956 0.74 1.156 0.812 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.284 0.412 1.44 0.484 ; 
RECT 1.368 0.412 1.44 0.812 ; 
RECT 1.368 0.74 1.532 0.812 ; 
END 
END A2 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.8 0.412 1.872 0.972 ; 
RECT 1.8 0.9 1.964 0.972 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.468 0.252 1.656 0.324 ; 
RECT 1.584 0.252 1.656 0.668 ; 
END 
END B2 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.284 0.108 0.364 0.972 ; 
RECT 0.284 0.9 0.48 0.972 ; 
RECT 0.284 0.108 0.488 0.18 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.16 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.16 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.72 0.252 1.344 0.324 ; 
RECT 0.56 0.504 0.792 0.576 ; 
RECT 0.72 0.252 0.792 0.972 ; 
RECT 0.72 0.9 1.568 0.972 ; 
RECT 1.024 0.108 2 0.18 ; 
END 
END OA22x2_ASAP7_75t_R 

MACRO OAI21xp5_ASAP7_75t_R_v1 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN OAI21xp5_ASAP7_75t_R_v1 0 0 ; 
SIZE 1.08 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.116 0.252 0.292 0.324 ; 
RECT 0.22 0.252 0.292 0.972 ; 
RECT 0.12 0.9 0.292 0.972 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.424 0.576 0.812 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.716 0.424 0.788 0.684 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.396 0.252 1.008 0.324 ; 
RECT 0.936 0.252 1.008 0.972 ; 
RECT 0.592 0.9 1.008 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.08 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.08 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.168 0.108 0.696 0.18 ; 
END 
END OAI21xp5_ASAP7_75t_R_v1 

MACRO OAI21xp5_ASAP7_75t_R_v2 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN OAI21xp5_ASAP7_75t_R_v2 0 0 ; 
SIZE 1.08 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.392 0.252 0.576 0.324 ; 
RECT 0.504 0.252 0.576 0.684 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.116 0.252 0.292 0.324 ; 
RECT 0.22 0.252 0.292 0.812 ; 
RECT 0.12 0.74 0.292 0.812 ; 
END 
END A2 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.788 0.412 0.86 0.812 ; 
RECT 0.692 0.74 0.86 0.812 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.824 0.108 1.008 0.18 ; 
RECT 0.936 0.108 1.008 0.972 ; 
RECT 0.16 0.9 1.008 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.08 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.08 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.168 0.108 0.688 0.18 ; 
END 
END OAI21xp5_ASAP7_75t_R_v2 

MACRO OAI22xp5_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN -0.216 0 ; 
FOREIGN OAI22xp5_ASAP7_75t_R 0.864 0 ; 
SIZE 1.296 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.084 0.412 1.156 0.812 ; 
RECT 1.084 0.412 1.252 0.484 ; 
RECT 1.084 0.74 1.252 0.812 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.368 0.476 1.44 0.812 ; 
RECT 1.368 0.74 1.532 0.812 ; 
END 
END A2 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.8 0.412 1.872 0.972 ; 
RECT 1.8 0.9 1.964 0.972 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.468 0.252 1.656 0.324 ; 
RECT 1.584 0.252 1.656 0.668 ; 
END 
END B2 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.94 0.252 1.012 0.972 ; 
RECT 0.94 0.252 1.344 0.324 ; 
RECT 0.94 0.9 1.568 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0.864 1.044 2.16 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0.864 -0.009 2.16 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 1.024 0.108 2 0.18 ; 
END 
END OAI22xp5_ASAP7_75t_R 

MACRO OAI31xp67_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN OAI31xp67_ASAP7_75t_R 0 0 ; 
SIZE 2.808 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.2 0.504 2.596 0.576 ; 
RECT 2.524 0.504 2.596 0.792 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.288 0.504 1.36 0.792 ; 
RECT 1.288 0.504 1.712 0.576 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.196 0.264 0.36 0.336 ; 
RECT 0.288 0.264 0.36 0.808 ; 
RECT 0.196 0.736 0.36 0.808 ; 
END 
END A3 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.624 0.284 0.696 0.8 ; 
RECT 0.624 0.504 0.852 0.576 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.104 0.9 2.688 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.808 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.808 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.384 0.9 1.788 0.972 ; 
RECT 0.164 0.108 2.216 0.18 ; 
RECT 1.464 0.696 2.424 0.768 ; 
RECT 2.484 0.108 2.704 0.18 ; 
RECT 2.632 0.108 2.704 0.36 ; 
RECT 0.796 0.288 2.704 0.36 ; 
RECT 1.04 0.288 1.112 0.828 ; 
RECT 0.8 0.756 1.112 0.828 ; 
END 
END OAI31xp67_ASAP7_75t_R 

MACRO OAI32xp33_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN OAI32xp33_ASAP7_75t_R 0 0 ; 
SIZE 1.728 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.132 0.108 0.292 0.18 ; 
RECT 0.22 0.108 0.292 0.828 ; 
RECT 0.132 0.756 0.292 0.828 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.416 0.268 0.576 0.352 ; 
RECT 0.504 0.268 0.576 0.828 ; 
RECT 0.416 0.756 0.576 0.828 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.268 0.792 0.672 ; 
RECT 0.72 0.268 0.888 0.34 ; 
END 
END A3 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.472 1.008 0.812 ; 
RECT 0.936 0.74 1.104 0.812 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.22 0.412 1.292 0.812 ; 
RECT 1.22 0.74 1.408 0.812 ; 
RECT 1.22 0.412 1.42 0.484 ; 
END 
END B2 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.04 0.252 1.604 0.324 ; 
RECT 1.532 0.252 1.604 0.972 ; 
RECT 0.16 0.9 1.604 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.728 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.728 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.392 0.108 1.336 0.18 ; 
END 
END OAI32xp33_ASAP7_75t_R 

MACRO OAI33xp33_ASAP_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN OAI33xp33_ASAP_75t_R 0 0 ; 
SIZE 1.944 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.068 0.504 0.14 0.972 ; 
RECT 0.068 0.9 0.252 0.972 ; 
RECT 0.068 0.504 0.36 0.576 ; 
RECT 0.288 0.504 0.36 0.648 ; 
END 
END A1 
PIN A2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.068 0.108 0.14 0.432 ; 
RECT 0.068 0.108 0.244 0.18 ; 
RECT 0.068 0.36 0.576 0.432 ; 
RECT 0.504 0.36 0.576 0.612 ; 
END 
END A2 
PIN A3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.72 0.252 0.792 0.6 ; 
RECT 0.72 0.252 0.892 0.324 ; 
END 
END A3 
PIN B1 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.936 0.516 1.008 0.812 ; 
RECT 0.832 0.736 1.008 0.812 ; 
END 
END B1 
PIN B2 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.152 0.5 1.224 0.812 ; 
RECT 1.152 0.74 1.328 0.812 ; 
END 
END B2 
PIN B3 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.436 0.4 1.508 0.668 ; 
RECT 1.436 0.4 1.608 0.472 ; 
RECT 1.436 0.596 1.608 0.668 ; 
END 
END B3 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.024 0.252 1.872 0.324 ; 
RECT 1.8 0.252 1.872 0.972 ; 
RECT 0.804 0.9 1.872 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.944 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.944 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.388 0.108 1.352 0.18 ; 
END 
END OAI33xp33_ASAP_75t_R 

MACRO SDFHx1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN SDFHx1_ASAP7_75t_R 0 0 ; 
SIZE 5.4 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.288 0.332 0.792 ; 
RECT 0.26 0.72 0.48 0.792 ; 
RECT 0.408 0.72 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.36 ; 
RECT 0.26 0.288 0.492 0.36 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.584 0.432 1.656 0.652 ; 
RECT 1.584 0.432 1.748 0.504 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 5.128 0.144 5.332 0.216 ; 
RECT 5.26 0.144 5.332 0.936 ; 
RECT 5.128 0.864 5.332 0.936 ; 
END 
END QN 
PIN SE 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M2 ; 
RECT 0.896 0.144 4.98 0.216 ; 
LAYER M1 ; 
RECT 0.868 0.144 0.94 0.576 ; 
RECT 0.868 0.144 1.032 0.216 ; 
RECT 0.868 0.504 1.192 0.576 ; 
RECT 4.824 0.144 4.896 0.668 ; 
RECT 4.824 0.144 5 0.216 ; 
LAYER V1 ; 
RECT 0.94 0.144 1.012 0.216 ; 
RECT 4.908 0.144 4.98 0.216 ; 
END 
END SE 
PIN SI 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.864 0.48 1.936 0.668 ; 
END 
END SI 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 5.4 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 5.4 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 1.368 0.288 1.532 0.36 ; 
RECT 1.368 0.288 1.44 0.596 ; 
RECT 1.236 0.752 1.788 0.824 ; 
RECT 1.02 0.9 2 0.972 ; 
RECT 1.16 0.108 2 0.18 ; 
RECT 1.16 0.108 1.232 0.384 ; 
RECT 1.04 0.312 1.232 0.384 ; 
RECT 2.104 0.504 2.332 0.576 ; 
RECT 2.104 0.504 2.216 0.792 ; 
RECT 1.668 0.28 2.436 0.352 ; 
RECT 2.448 0.44 2.52 0.696 ; 
RECT 2.88 0.66 2.952 0.812 ; 
RECT 2.536 0.108 2.736 0.18 ; 
RECT 2.664 0.488 3.176 0.56 ; 
RECT 2.664 0.108 2.736 0.956 ; 
RECT 2.32 0.884 2.736 0.956 ; 
RECT 3.204 0.18 3.276 0.416 ; 
RECT 2.848 0.344 3.408 0.416 ; 
RECT 3.336 0.344 3.408 0.968 ; 
RECT 3.168 0.896 3.408 0.968 ; 
RECT 3.528 0.404 3.6 0.668 ; 
RECT 3.4 0.108 3.816 0.18 ; 
RECT 4.176 0.468 4.248 0.692 ; 
RECT 3.744 0.62 4.248 0.692 ; 
RECT 3.744 0.108 3.816 0.968 ; 
RECT 3.616 0.896 3.816 0.968 ; 
RECT 3.96 0.108 4.464 0.18 ; 
RECT 3.96 0.108 4.032 0.476 ; 
RECT 4.392 0.108 4.464 0.968 ; 
RECT 4.264 0.896 4.464 0.968 ; 
RECT 4.604 0.136 4.676 0.972 ; 
RECT 4.604 0.9 4.808 0.972 ; 
RECT 5.04 0.36 5.112 0.668 ; 
LAYER M2 ; 
RECT 0.704 0.72 2.952 0.792 ; 
RECT 0.076 0.576 3.6 0.648 ; 
RECT 1.396 0.288 4.676 0.36 ; 
RECT 3.744 0.576 5.132 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 0.94 0.144 1.012 0.216 ; 
RECT 1.44 0.288 1.512 0.36 ; 
RECT 2.124 0.72 2.196 0.792 ; 
RECT 2.448 0.576 2.52 0.648 ; 
RECT 2.88 0.72 2.952 0.792 ; 
RECT 3.528 0.576 3.6 0.648 ; 
RECT 3.744 0.576 3.816 0.648 ; 
RECT 4.604 0.288 4.676 0.36 ; 
RECT 4.908 0.144 4.98 0.216 ; 
RECT 5.04 0.576 5.112 0.648 ; 
END 
END SDFHx1_ASAP7_75t_R 

MACRO SDFHx3_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN SDFHx3_ASAP7_75t_R 0 0 ; 
SIZE 6.912 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.26 0.288 0.332 0.792 ; 
RECT 0.26 0.72 0.48 0.792 ; 
RECT 0.408 0.72 0.48 0.944 ; 
RECT 0.42 0.14 0.492 0.36 ; 
RECT 0.26 0.288 0.492 0.36 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.78 0.576 1.852 0.936 ; 
RECT 1.78 0.864 1.984 0.936 ; 
RECT 1.952 0.464 2.024 0.648 ; 
RECT 1.78 0.576 2.024 0.648 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 6.204 0.144 6.844 0.216 ; 
RECT 6.772 0.144 6.844 0.936 ; 
RECT 6.204 0.864 6.844 0.936 ; 
END 
END QN 
PIN SE 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.124 0.288 1.196 0.792 ; 
RECT 1.124 0.72 1.344 0.792 ; 
RECT 1.272 0.72 1.344 0.944 ; 
RECT 1.284 0.14 1.356 0.36 ; 
RECT 1.124 0.288 1.356 0.36 ; 
END 
END SE 
PIN SI 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 3.096 0.288 3.168 0.628 ; 
RECT 3.56 0.14 3.632 0.36 ; 
RECT 3.096 0.288 3.632 0.36 ; 
END 
END SI 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 6.912 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 6.912 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.076 0.108 0.272 0.18 ; 
RECT 0.076 0.108 0.148 0.972 ; 
RECT 0.076 0.9 0.272 0.972 ; 
RECT 0.568 0.488 0.64 0.668 ; 
RECT 0.592 0.108 0.796 0.18 ; 
RECT 0.724 0.108 0.796 0.972 ; 
RECT 0.592 0.9 0.796 0.972 ; 
RECT 0.94 0.108 1.136 0.18 ; 
RECT 0.94 0.108 1.012 0.972 ; 
RECT 0.94 0.9 1.136 0.972 ; 
RECT 1.432 0.412 1.504 0.652 ; 
RECT 1.456 0.108 1.66 0.18 ; 
RECT 1.588 0.108 1.66 0.972 ; 
RECT 1.456 0.9 1.66 0.972 ; 
RECT 2.3 0.412 2.372 0.58 ; 
RECT 2.208 0.508 2.372 0.58 ; 
RECT 2.472 0.288 2.76 0.36 ; 
RECT 2.548 0.288 2.62 0.572 ; 
RECT 2.548 0.5 2.992 0.572 ; 
RECT 2.104 0.72 3.08 0.792 ; 
RECT 2.752 0.9 3.296 0.972 ; 
RECT 1.888 0.112 3.296 0.184 ; 
RECT 3.528 0.468 3.6 0.812 ; 
RECT 3.744 0.432 3.816 0.668 ; 
RECT 4.176 0.66 4.248 0.812 ; 
RECT 3.832 0.108 4.032 0.18 ; 
RECT 3.96 0.488 4.472 0.56 ; 
RECT 3.96 0.108 4.032 0.972 ; 
RECT 3.616 0.9 4.032 0.972 ; 
RECT 4.5 0.18 4.572 0.416 ; 
RECT 4.144 0.344 4.704 0.416 ; 
RECT 4.632 0.344 4.704 0.968 ; 
RECT 4.464 0.896 4.704 0.968 ; 
RECT 4.824 0.404 4.896 0.668 ; 
RECT 4.696 0.108 5.112 0.18 ; 
RECT 5.472 0.468 5.544 0.692 ; 
RECT 5.04 0.62 5.544 0.692 ; 
RECT 5.04 0.108 5.112 0.968 ; 
RECT 4.912 0.896 5.112 0.968 ; 
RECT 5.256 0.108 5.76 0.18 ; 
RECT 5.256 0.108 5.328 0.476 ; 
RECT 5.688 0.108 5.76 0.968 ; 
RECT 5.56 0.896 5.76 0.968 ; 
RECT 6.12 0.36 6.192 0.668 ; 
LAYER M2 ; 
RECT 0.932 0.432 2.4 0.504 ; 
RECT 1.572 0.288 2.64 0.36 ; 
RECT 0.712 0.72 4.268 0.792 ; 
RECT 0.064 0.576 4.896 0.648 ; 
RECT 5.04 0.576 6.212 0.648 ; 
LAYER V1 ; 
RECT 0.076 0.576 0.148 0.648 ; 
RECT 0.568 0.576 0.64 0.648 ; 
RECT 0.724 0.72 0.796 0.792 ; 
RECT 0.94 0.432 1.012 0.504 ; 
RECT 1.432 0.432 1.504 0.504 ; 
RECT 1.588 0.288 1.66 0.36 ; 
RECT 2.3 0.432 2.372 0.504 ; 
RECT 2.548 0.288 2.62 0.36 ; 
RECT 3.528 0.72 3.6 0.792 ; 
RECT 3.744 0.576 3.816 0.648 ; 
RECT 4.176 0.72 4.248 0.792 ; 
RECT 4.824 0.576 4.896 0.648 ; 
RECT 5.04 0.576 5.112 0.648 ; 
RECT 6.12 0.576 6.192 0.648 ; 
END 
END SDFHx3_ASAP7_75t_R 

MACRO SDFHx4_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN SDFHx4_ASAP7_75t_R 0 0 ; 
SIZE 6.912 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.452 0.36 0.716 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.512 0.432 1.584 0.936 ; 
RECT 1.512 0.432 1.872 0.504 ; 
RECT 1.512 0.864 1.836 0.936 ; 
RECT 1.8 0.432 1.872 0.596 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 5.776 0.144 6.804 0.216 ; 
RECT 6.732 0.144 6.804 0.936 ; 
RECT 5.776 0.864 6.804 0.936 ; 
END 
END QN 
PIN SE 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M2 ; 
RECT 0.86 0.288 2.5 0.36 ; 
LAYER M1 ; 
RECT 0.856 0.144 1.024 0.216 ; 
RECT 0.952 0.144 1.024 0.36 ; 
RECT 0.952 0.288 1.156 0.36 ; 
RECT 1.084 0.288 1.156 0.936 ; 
RECT 0.948 0.864 1.156 0.936 ; 
RECT 2.232 0.288 2.304 0.596 ; 
RECT 2.232 0.288 2.396 0.36 ; 
LAYER V1 ; 
RECT 1.012 0.288 1.084 0.36 ; 
RECT 2.304 0.288 2.376 0.36 ; 
END 
END SE 
PIN SI 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.448 0.432 2.52 0.596 ; 
RECT 2.56 0.288 2.632 0.504 ; 
RECT 2.448 0.432 2.632 0.504 ; 
RECT 2.78 0.144 2.852 0.36 ; 
RECT 2.56 0.288 2.852 0.36 ; 
RECT 2.78 0.144 3.068 0.216 ; 
END 
END SI 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 6.912 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 6.912 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.108 0.108 0.34 0.18 ; 
RECT 0.268 0.108 0.34 0.336 ; 
RECT 0.268 0.264 0.576 0.336 ; 
RECT 0.504 0.264 0.576 0.716 ; 
RECT 0.108 0.108 0.18 0.972 ; 
RECT 0.108 0.9 0.272 0.972 ; 
RECT 0.592 0.108 0.756 0.18 ; 
RECT 0.684 0.108 0.756 0.972 ; 
RECT 0.592 0.9 0.756 0.972 ; 
RECT 1.26 0.288 2.088 0.36 ; 
RECT 2.016 0.288 2.088 0.596 ; 
RECT 1.26 0.18 1.332 0.88 ; 
RECT 1.684 0.696 2.648 0.768 ; 
RECT 1.672 0.108 2.648 0.18 ; 
RECT 2.732 0.484 2.804 0.668 ; 
RECT 2.32 0.9 3.08 0.972 ; 
RECT 3.096 0.408 3.168 0.596 ; 
RECT 3.312 0.484 3.384 0.668 ; 
RECT 2.952 0.34 3.024 0.828 ; 
RECT 2.952 0.756 3.276 0.828 ; 
RECT 3.204 0.756 3.276 0.972 ; 
RECT 3.744 0.484 3.816 0.972 ; 
RECT 3.204 0.9 3.816 0.972 ; 
RECT 3.528 0.256 4.036 0.328 ; 
RECT 3.528 0.256 3.6 0.596 ; 
RECT 3.964 0.256 4.036 0.916 ; 
RECT 4.392 0.484 4.464 0.672 ; 
RECT 4.608 0.408 4.68 0.596 ; 
RECT 4.824 0.484 4.896 0.672 ; 
RECT 5.04 0.484 5.112 0.968 ; 
RECT 5.436 0.34 5.508 0.968 ; 
RECT 5.04 0.896 5.508 0.968 ; 
RECT 4.176 0.108 5.676 0.18 ; 
RECT 5.604 0.108 5.676 0.364 ; 
RECT 5.604 0.292 5.908 0.364 ; 
RECT 5.256 0.108 5.328 0.596 ; 
RECT 5.836 0.292 5.908 0.716 ; 
RECT 4.176 0.108 4.248 0.972 ; 
RECT 4.176 0.9 4.592 0.972 ; 
LAYER M2 ; 
RECT 0.636 0.432 4.744 0.504 ; 
RECT 0.436 0.576 4.968 0.648 ; 
LAYER V1 ; 
RECT 0.504 0.576 0.576 0.648 ; 
RECT 0.684 0.432 0.756 0.504 ; 
RECT 1.012 0.288 1.084 0.36 ; 
RECT 2.304 0.288 2.376 0.36 ; 
RECT 2.732 0.576 2.804 0.648 ; 
RECT 3.096 0.432 3.168 0.504 ; 
RECT 3.312 0.576 3.384 0.648 ; 
RECT 4.392 0.576 4.464 0.648 ; 
RECT 4.608 0.432 4.68 0.504 ; 
RECT 4.824 0.576 4.896 0.648 ; 
END 
END SDFHx4_ASAP7_75t_R 

MACRO SDFLx1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN SDFLx1_ASAP7_75t_R 0 0 ; 
SIZE 6.48 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN CLK 
DIRECTION INPUT ; 
USE CLOCK ; 
PORT 
LAYER M1 ; 
RECT 2.852 0.388 2.924 0.648 ; 
RECT 2.852 0.576 3.016 0.648 ; 
END 
END CLK 
PIN D 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.88 0.472 0.952 0.792 ; 
RECT 0.748 0.72 0.952 0.792 ; 
END 
END D 
PIN QN 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 6.208 0.144 6.412 0.216 ; 
RECT 6.34 0.144 6.412 0.936 ; 
RECT 6.208 0.864 6.412 0.936 ; 
END 
END QN 
PIN SE 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M2 ; 
RECT 0.28 0.432 1.656 0.504 ; 
LAYER M1 ; 
RECT 0.072 0.144 0.144 0.416 ; 
RECT 0.072 0.144 0.252 0.216 ; 
RECT 0.072 0.344 0.36 0.416 ; 
RECT 0.288 0.344 0.36 0.792 ; 
RECT 0.108 0.72 0.36 0.792 ; 
RECT 1.584 0.412 1.656 0.596 ; 
LAYER V1 ; 
RECT 0.288 0.432 0.36 0.504 ; 
RECT 1.584 0.432 1.656 0.504 ; 
END 
END SE 
PIN SI 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.372 0.252 1.444 0.604 ; 
RECT 1.372 0.252 1.56 0.324 ; 
END 
END SI 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 6.48 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 6.48 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.376 0.108 0.576 0.18 ; 
RECT 0.504 0.26 1.224 0.332 ; 
RECT 1.152 0.26 1.224 0.648 ; 
RECT 0.504 0.108 0.576 0.972 ; 
RECT 0.376 0.9 0.576 0.972 ; 
RECT 0.816 0.108 1.768 0.18 ; 
RECT 0.816 0.896 1.776 0.968 ; 
RECT 1.8 0.412 1.872 0.592 ; 
RECT 1.464 0.744 2.208 0.816 ; 
RECT 2.236 0.476 2.308 0.668 ; 
RECT 1.908 0.204 2.524 0.276 ; 
RECT 2.452 0.204 2.524 0.936 ; 
RECT 2.324 0.864 2.524 0.936 ; 
RECT 2.668 0.108 2.864 0.18 ; 
RECT 3.16 0.488 3.232 0.792 ; 
RECT 2.668 0.72 3.232 0.792 ; 
RECT 2.668 0.108 2.74 0.972 ; 
RECT 2.668 0.9 2.864 0.972 ; 
RECT 3.184 0.108 3.388 0.18 ; 
RECT 3.316 0.432 3.816 0.504 ; 
RECT 3.744 0.432 3.816 0.668 ; 
RECT 3.316 0.108 3.388 0.972 ; 
RECT 3.184 0.9 3.388 0.972 ; 
RECT 4.176 0.66 4.248 0.812 ; 
RECT 3.832 0.108 4.032 0.18 ; 
RECT 3.96 0.488 4.472 0.56 ; 
RECT 3.96 0.108 4.032 0.936 ; 
RECT 3.524 0.864 4.032 0.936 ; 
RECT 4.5 0.18 4.572 0.416 ; 
RECT 4.144 0.344 4.704 0.416 ; 
RECT 4.632 0.344 4.704 0.968 ; 
RECT 4.464 0.896 4.704 0.968 ; 
RECT 4.824 0.436 4.896 0.7 ; 
RECT 4.696 0.108 5.112 0.18 ; 
RECT 5.472 0.468 5.544 0.692 ; 
RECT 5.04 0.62 5.544 0.692 ; 
RECT 5.04 0.108 5.112 0.968 ; 
RECT 4.912 0.896 5.112 0.968 ; 
RECT 5.256 0.108 5.76 0.18 ; 
RECT 5.256 0.108 5.328 0.476 ; 
RECT 5.688 0.108 5.76 0.968 ; 
RECT 5.56 0.896 5.76 0.968 ; 
RECT 6.12 0.36 6.192 0.668 ; 
LAYER M2 ; 
RECT 2.228 0.576 2.744 0.648 ; 
RECT 1.8 0.432 3.392 0.504 ; 
RECT 2.424 0.864 3.632 0.936 ; 
RECT 2.452 0.288 4.032 0.36 ; 
RECT 3.068 0.72 4.252 0.792 ; 
RECT 3.716 0.576 4.912 0.648 ; 
RECT 5.04 0.576 6.204 0.648 ; 
LAYER V1 ; 
RECT 0.288 0.432 0.36 0.504 ; 
RECT 1.584 0.432 1.656 0.504 ; 
RECT 1.8 0.432 1.872 0.504 ; 
RECT 2.236 0.576 2.308 0.648 ; 
RECT 2.424 0.864 2.496 0.936 ; 
RECT 2.452 0.288 2.524 0.36 ; 
RECT 2.668 0.576 2.74 0.648 ; 
RECT 3.076 0.72 3.148 0.792 ; 
RECT 3.316 0.432 3.388 0.504 ; 
RECT 3.548 0.864 3.62 0.936 ; 
RECT 3.744 0.576 3.816 0.648 ; 
RECT 3.96 0.288 4.032 0.36 ; 
RECT 4.176 0.72 4.248 0.792 ; 
RECT 4.824 0.576 4.896 0.648 ; 
RECT 5.04 0.576 5.112 0.648 ; 
RECT 6.12 0.576 6.192 0.648 ; 
END 
END SDFLx1_ASAP7_75t_R 

MACRO TAPCELL_ASAP7_75t 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN TAPCELL_ASAP7_75t 0 0 ; 
SIZE 0.432 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 0.432 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 0.432 0.036 ; 
END 
END vss! 
END TAPCELL_ASAP7_75t 

MACRO XNOR2xp5_ASAP7_75t_R_v1 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN XNOR2xp5_ASAP7_75t_R_v1 0 0 ; 
SIZE 3.024 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.288 0.252 0.36 0.772 ; 
RECT 0.288 0.7 0.684 0.772 ; 
RECT 0.612 0.7 0.684 0.972 ; 
RECT 0.612 0.9 0.792 0.972 ; 
RECT 0.288 0.252 0.9 0.324 ; 
RECT 0.828 0.252 0.9 0.58 ; 
RECT 0.828 0.508 1.224 0.58 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.384 0.5 2.456 0.972 ; 
RECT 2.384 0.9 2.58 0.972 ; 
RECT 2.564 0.288 2.64 0.572 ; 
RECT 2.564 0.288 2.748 0.36 ; 
RECT 2.384 0.5 2.748 0.572 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.04 0.256 1.552 0.328 ; 
RECT 1.48 0.256 1.552 0.828 ; 
RECT 1.26 0.756 1.764 0.828 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 3.024 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 3.024 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.072 0.108 0.692 0.18 ; 
RECT 0.072 0.108 0.144 0.972 ; 
RECT 0.072 0.9 0.284 0.972 ; 
RECT 1.04 0.9 1.984 0.972 ; 
RECT 0.82 0.108 2.212 0.18 ; 
RECT 2.376 0.108 2.948 0.18 ; 
RECT 2.376 0.108 2.448 0.324 ; 
RECT 1.8 0.252 2.448 0.324 ; 
RECT 1.8 0.252 1.872 0.596 ; 
RECT 2.876 0.108 2.948 0.796 ; 
RECT 2.748 0.724 2.948 0.796 ; 
END 
END XNOR2xp5_ASAP7_75t_R_v1 

MACRO XNOR2xp5_ASAP7_75t_R_v2 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN XNOR2xp5_ASAP7_75t_R_v2 0 0 ; 
SIZE 1.944 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.22 0.108 0.292 0.812 ; 
RECT 0.116 0.74 0.292 0.812 ; 
RECT 0.22 0.108 0.884 0.18 ; 
RECT 0.812 0.108 0.884 0.324 ; 
RECT 0.812 0.252 1.44 0.324 ; 
RECT 1.368 0.252 1.44 0.6 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.424 0.268 0.576 0.34 ; 
RECT 0.504 0.268 0.576 0.812 ; 
RECT 0.428 0.74 0.576 0.812 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.688 0.108 1.872 0.18 ; 
RECT 1.8 0.108 1.872 0.972 ; 
RECT 1.024 0.9 1.872 0.972 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 1.944 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 1.944 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 1.04 0.108 1.552 0.18 ; 
RECT 1.652 0.488 1.724 0.812 ; 
RECT 0.648 0.74 1.724 0.812 ; 
RECT 0.648 0.332 0.72 0.972 ; 
RECT 0.376 0.9 0.72 0.972 ; 
END 
END XNOR2xp5_ASAP7_75t_R_v2 

MACRO XOR2x1_ASAP7_75t_R 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN XOR2x1_ASAP7_75t_R 0 0 ; 
SIZE 4.104 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.224 0.256 0.296 0.792 ; 
RECT 1.156 0.492 1.228 0.792 ; 
RECT 0.224 0.72 1.228 0.792 ; 
RECT 1.156 0.588 1.888 0.66 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.504 0.484 0.576 0.648 ; 
RECT 1.008 0.288 1.08 0.648 ; 
RECT 0.504 0.576 1.08 0.648 ; 
RECT 1.008 0.288 1.66 0.36 ; 
RECT 1.588 0.288 1.66 0.476 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.592 0.108 4.032 0.18 ; 
RECT 3.96 0.108 4.032 0.788 ; 
RECT 3.184 0.716 4.032 0.788 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 4.104 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 4.104 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.396 0.252 0.908 0.324 ; 
RECT 0.396 0.252 0.468 0.4 ; 
RECT 2.876 0.664 2.948 0.828 ; 
RECT 1.384 0.756 2.948 0.828 ; 
RECT 2.536 0.292 3.728 0.364 ; 
RECT 1.888 0.252 2.232 0.324 ; 
RECT 2.16 0.492 3.82 0.564 ; 
RECT 2.16 0.252 2.232 0.66 ; 
RECT 2.028 0.588 2.232 0.66 ; 
RECT 0.16 0.9 3.944 0.972 ; 
END 
END XOR2x1_ASAP7_75t_R 

MACRO XOR2xp5_ASAP7_75t_R_v1 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN XOR2xp5_ASAP7_75t_R_v1 0 0 ; 
SIZE 2.808 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.18 0.268 0.252 0.832 ; 
RECT 0.18 0.504 1.244 0.576 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.564 0.504 2.628 0.576 ; 
RECT 2.556 0.288 2.628 0.832 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.024 0.308 1.44 0.38 ; 
RECT 1.368 0.308 1.44 0.812 ; 
RECT 1.24 0.74 1.44 0.812 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.808 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.808 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 1.032 0.9 1.772 0.972 ; 
RECT 0.808 0.108 2 0.18 ; 
END 
END XOR2xp5_ASAP7_75t_R_v1 

MACRO XOR2xp5_ASAP7_75t_R_v2 
CLASS CORE ; 
ORIGIN 0 0 ; 
FOREIGN XOR2xp5_ASAP7_75t_R_v2 0 0 ; 
SIZE 2.808 BY 1.08 ; 
SYMMETRY X Y ; 
SITE coreSite ; 
PIN A 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 0.368 0.288 0.44 0.792 ; 
RECT 0.272 0.72 0.44 0.792 ; 
RECT 0.368 0.288 0.58 0.36 ; 
RECT 0.268 0.504 1.02 0.576 ; 
END 
END A 
PIN B 
DIRECTION INPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 2.34 0.288 2.412 0.792 ; 
RECT 2.2 0.72 2.412 0.792 ; 
RECT 2.34 0.288 2.516 0.36 ; 
RECT 1.788 0.504 2.54 0.576 ; 
END 
END B 
PIN Y 
DIRECTION OUTPUT ; 
USE SIGNAL ; 
PORT 
LAYER M1 ; 
RECT 1.016 0.288 1.44 0.36 ; 
RECT 1.368 0.288 1.44 0.792 ; 
RECT 1.368 0.72 1.568 0.792 ; 
END 
END Y 
PIN vdd! 
DIRECTION INOUT ; 
USE POWER ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 1.044 2.808 1.116 ; 
END 
END vdd! 
PIN vss! 
DIRECTION INOUT ; 
USE GROUND ; 
SHAPE ABUTMENT ; 
PORT 
LAYER M1 ; 
RECT 0 -0.009 2.808 0.036 ; 
END 
END vss! 
OBS 
LAYER M1 ; 
RECT 0.072 0.108 0.268 0.18 ; 
RECT 1.152 0.484 1.224 0.828 ; 
RECT 0.72 0.756 1.224 0.828 ; 
RECT 0.072 0.108 0.144 0.972 ; 
RECT 0.72 0.756 0.792 0.972 ; 
RECT 0.072 0.9 0.792 0.972 ; 
RECT 1.02 0.9 1.784 0.972 ; 
RECT 0.804 0.108 2 0.18 ; 
RECT 2.132 0.108 2.736 0.18 ; 
RECT 2.132 0.108 2.204 0.324 ; 
RECT 1.584 0.252 2.204 0.324 ; 
RECT 1.584 0.252 1.656 0.592 ; 
RECT 2.664 0.108 2.736 0.972 ; 
RECT 2.536 0.9 2.736 0.972 ; 
END 
END XOR2xp5_ASAP7_75t_R_v2 

END LIBRARY 
